<?xml version="1.0" encoding="UTF-8"?>
<svg xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" width="504pt" height="504pt" viewBox="0 0 504 504" version="1.1">
<defs>
<g>
<symbol overflow="visible" id="glyph0-0">
<path style="stroke:none;" d="M 1.800781 0 L 1.800781 -9 L 9 -9 L 9 0 Z M 2.023438 -0.226563 L 8.773438 -0.226563 L 8.773438 -8.773438 L 2.023438 -8.773438 Z M 2.023438 -0.226563 "/>
</symbol>
<symbol overflow="visible" id="glyph0-1">
<path style="stroke:none;" d="M 1.070313 0 L 1.070313 -10.308594 L 3.09375 -10.308594 L 7.3125 -3.425781 L 7.3125 -10.308594 L 9.246094 -10.308594 L 9.246094 0 L 7.15625 0 L 3.003906 -6.722656 L 3.003906 0 Z M 1.070313 0 "/>
</symbol>
<symbol overflow="visible" id="glyph0-2">
<path style="stroke:none;" d="M 5.949219 0 L 5.949219 -1.117188 C 5.671875 -0.714844 5.316406 -0.402344 4.875 -0.175781 C 4.429688 0.0507813 3.960938 0.164063 3.472656 0.167969 C 2.96875 0.164063 2.519531 0.0585938 2.125 -0.160156 C 1.722656 -0.378906 1.433594 -0.691406 1.257813 -1.089844 C 1.078125 -1.488281 0.988281 -2.039063 0.992188 -2.742188 L 0.992188 -7.46875 L 2.96875 -7.46875 L 2.96875 -4.035156 C 2.964844 -2.984375 3 -2.339844 3.074219 -2.105469 C 3.144531 -1.863281 3.277344 -1.675781 3.472656 -1.542969 C 3.664063 -1.402344 3.90625 -1.335938 4.203125 -1.335938 C 4.539063 -1.335938 4.84375 -1.425781 5.109375 -1.613281 C 5.375 -1.792969 5.558594 -2.023438 5.660156 -2.300781 C 5.757813 -2.574219 5.804688 -3.246094 5.808594 -4.316406 L 5.808594 -7.46875 L 7.785156 -7.46875 L 7.785156 0 Z M 5.949219 0 "/>
</symbol>
<symbol overflow="visible" id="glyph0-3">
<path style="stroke:none;" d="M 0.886719 -7.46875 L 2.707031 -7.46875 L 2.707031 -6.449219 C 3.355469 -7.238281 4.128906 -7.632813 5.035156 -7.636719 C 5.507813 -7.632813 5.921875 -7.535156 6.277344 -7.339844 C 6.625 -7.140625 6.914063 -6.84375 7.144531 -6.449219 C 7.46875 -6.84375 7.824219 -7.140625 8.203125 -7.339844 C 8.582031 -7.535156 8.988281 -7.632813 9.421875 -7.636719 C 9.96875 -7.632813 10.429688 -7.523438 10.8125 -7.300781 C 11.1875 -7.078125 11.472656 -6.75 11.664063 -6.320313 C 11.796875 -6 11.863281 -5.484375 11.867188 -4.773438 L 11.867188 0 L 9.894531 0 L 9.894531 -4.269531 C 9.890625 -5.007813 9.820313 -5.484375 9.6875 -5.703125 C 9.5 -5.980469 9.21875 -6.121094 8.84375 -6.125 C 8.5625 -6.121094 8.304688 -6.039063 8.0625 -5.871094 C 7.820313 -5.699219 7.644531 -5.449219 7.535156 -5.128906 C 7.425781 -4.800781 7.371094 -4.289063 7.375 -3.585938 L 7.375 0 L 5.398438 0 L 5.398438 -4.09375 C 5.394531 -4.816406 5.359375 -5.285156 5.292969 -5.5 C 5.21875 -5.707031 5.109375 -5.863281 4.964844 -5.96875 C 4.816406 -6.070313 4.617188 -6.121094 4.367188 -6.125 C 4.058594 -6.121094 3.785156 -6.039063 3.542969 -5.878906 C 3.296875 -5.710938 3.121094 -5.476563 3.019531 -5.167969 C 2.910156 -4.855469 2.859375 -4.339844 2.863281 -3.628906 L 2.863281 0 L 0.886719 0 Z M 0.886719 -7.46875 "/>
</symbol>
<symbol overflow="visible" id="glyph1-0">
<path style="stroke:none;" d="M 1.5 0 L 1.5 -7.5 L 7.5 -7.5 L 7.5 0 Z M 1.6875 -0.1875 L 7.3125 -0.1875 L 7.3125 -7.3125 L 1.6875 -7.3125 Z M 1.6875 -0.1875 "/>
</symbol>
<symbol overflow="visible" id="glyph1-1">
<path style="stroke:none;" d="M -0.015625 0 L 3.28125 -8.589844 L 4.507813 -8.589844 L 8.023438 0 L 6.726563 0 L 5.726563 -2.601563 L 2.132813 -2.601563 L 1.1875 0 Z M 2.460938 -3.527344 L 5.375 -3.527344 L 4.476563 -5.90625 C 4.203125 -6.628906 4 -7.222656 3.867188 -7.6875 C 3.757813 -7.132813 3.601563 -6.585938 3.40625 -6.046875 Z M 2.460938 -3.527344 "/>
</symbol>
<symbol overflow="visible" id="glyph1-2">
<path style="stroke:none;" d="M 2.519531 0 L 0.152344 -6.222656 L 1.265625 -6.222656 L 2.601563 -2.496094 C 2.746094 -2.089844 2.878906 -1.671875 3 -1.242188 C 3.09375 -1.570313 3.222656 -1.964844 3.390625 -2.425781 L 4.773438 -6.222656 L 5.859375 -6.222656 L 3.503906 0 Z M 2.519531 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-3">
<path style="stroke:none;" d="M 5.050781 -2.003906 L 6.140625 -1.867188 C 5.96875 -1.230469 5.648438 -0.738281 5.183594 -0.386719 C 4.71875 -0.0351563 4.125 0.140625 3.40625 0.140625 C 2.492188 0.140625 1.769531 -0.136719 1.238281 -0.699219 C 0.699219 -1.253906 0.433594 -2.042969 0.4375 -3.058594 C 0.433594 -4.105469 0.703125 -4.917969 1.246094 -5.496094 C 1.78125 -6.074219 2.480469 -6.363281 3.34375 -6.363281 C 4.175781 -6.363281 4.855469 -6.078125 5.382813 -5.511719 C 5.910156 -4.945313 6.175781 -4.148438 6.175781 -3.125 C 6.175781 -3.058594 6.171875 -2.964844 6.171875 -2.84375 L 1.53125 -2.84375 C 1.5625 -2.15625 1.757813 -1.632813 2.109375 -1.269531 C 2.457031 -0.90625 2.890625 -0.726563 3.410156 -0.726563 C 3.796875 -0.726563 4.125 -0.828125 4.402344 -1.03125 C 4.671875 -1.234375 4.890625 -1.558594 5.050781 -2.003906 Z M 1.585938 -3.710938 L 5.0625 -3.710938 C 5.015625 -4.226563 4.882813 -4.621094 4.664063 -4.886719 C 4.328125 -5.292969 3.890625 -5.496094 3.359375 -5.496094 C 2.871094 -5.496094 2.464844 -5.332031 2.136719 -5.007813 C 1.804688 -4.683594 1.621094 -4.25 1.585938 -3.710938 Z M 1.585938 -3.710938 "/>
</symbol>
<symbol overflow="visible" id="glyph1-4">
<path style="stroke:none;" d="M 0.78125 0 L 0.78125 -6.222656 L 1.726563 -6.222656 L 1.726563 -5.28125 C 1.96875 -5.71875 2.191406 -6.011719 2.398438 -6.152344 C 2.601563 -6.292969 2.828125 -6.363281 3.078125 -6.363281 C 3.429688 -6.363281 3.792969 -6.25 4.160156 -6.023438 L 3.796875 -5.046875 C 3.539063 -5.195313 3.28125 -5.273438 3.023438 -5.273438 C 2.792969 -5.273438 2.585938 -5.203125 2.402344 -5.066406 C 2.214844 -4.925781 2.082031 -4.734375 2.007813 -4.488281 C 1.890625 -4.113281 1.832031 -3.703125 1.835938 -3.257813 L 1.835938 0 Z M 0.78125 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-5">
<path style="stroke:none;" d="M 4.851563 -0.765625 C 4.460938 -0.433594 4.082031 -0.199219 3.722656 -0.0625 C 3.355469 0.0742188 2.96875 0.140625 2.5625 0.140625 C 1.875 0.140625 1.351563 -0.0234375 0.984375 -0.359375 C 0.617188 -0.6875 0.433594 -1.117188 0.433594 -1.640625 C 0.433594 -1.945313 0.5 -2.222656 0.640625 -2.472656 C 0.777344 -2.722656 0.960938 -2.925781 1.1875 -3.082031 C 1.410156 -3.234375 1.664063 -3.347656 1.945313 -3.429688 C 2.152344 -3.476563 2.464844 -3.53125 2.882813 -3.585938 C 3.734375 -3.6875 4.359375 -3.808594 4.765625 -3.949219 C 4.765625 -4.089844 4.769531 -4.179688 4.769531 -4.226563 C 4.769531 -4.648438 4.667969 -4.953125 4.46875 -5.132813 C 4.199219 -5.371094 3.800781 -5.488281 3.269531 -5.492188 C 2.769531 -5.488281 2.402344 -5.402344 2.167969 -5.230469 C 1.933594 -5.054688 1.757813 -4.746094 1.648438 -4.304688 L 0.617188 -4.445313 C 0.707031 -4.886719 0.863281 -5.242188 1.078125 -5.515625 C 1.289063 -5.78125 1.597656 -5.992188 2.007813 -6.140625 C 2.410156 -6.289063 2.882813 -6.363281 3.421875 -6.363281 C 3.953125 -6.363281 4.382813 -6.300781 4.714844 -6.175781 C 5.046875 -6.050781 5.292969 -5.890625 5.449219 -5.703125 C 5.605469 -5.511719 5.714844 -5.273438 5.777344 -4.984375 C 5.808594 -4.804688 5.824219 -4.480469 5.828125 -4.015625 L 5.828125 -2.609375 C 5.824219 -1.625 5.847656 -1.003906 5.894531 -0.746094 C 5.941406 -0.484375 6.03125 -0.238281 6.164063 0 L 5.0625 0 C 4.953125 -0.21875 4.882813 -0.472656 4.851563 -0.765625 Z M 4.765625 -3.125 C 4.375 -2.964844 3.800781 -2.832031 3.039063 -2.726563 C 2.605469 -2.660156 2.300781 -2.589844 2.121094 -2.515625 C 1.941406 -2.433594 1.800781 -2.320313 1.703125 -2.171875 C 1.605469 -2.019531 1.558594 -1.851563 1.558594 -1.671875 C 1.558594 -1.386719 1.664063 -1.152344 1.875 -0.96875 C 2.085938 -0.777344 2.398438 -0.683594 2.8125 -0.6875 C 3.21875 -0.683594 3.578125 -0.773438 3.894531 -0.953125 C 4.210938 -1.128906 4.445313 -1.371094 4.59375 -1.679688 C 4.707031 -1.917969 4.761719 -2.269531 4.765625 -2.734375 Z M 4.765625 -3.125 "/>
</symbol>
<symbol overflow="visible" id="glyph1-6">
<path style="stroke:none;" d="M 0.597656 0.515625 L 1.625 0.667969 C 1.664063 0.980469 1.785156 1.210938 1.980469 1.359375 C 2.242188 1.554688 2.597656 1.652344 3.054688 1.652344 C 3.539063 1.652344 3.917969 1.554688 4.183594 1.359375 C 4.449219 1.164063 4.628906 0.890625 4.722656 0.539063 C 4.777344 0.324219 4.800781 -0.125 4.796875 -0.8125 C 4.335938 -0.269531 3.761719 0 3.078125 0 C 2.21875 0 1.558594 -0.308594 1.089844 -0.925781 C 0.621094 -1.542969 0.386719 -2.28125 0.386719 -3.148438 C 0.386719 -3.738281 0.492188 -4.285156 0.707031 -4.789063 C 0.921875 -5.289063 1.234375 -5.679688 1.644531 -5.953125 C 2.050781 -6.226563 2.53125 -6.363281 3.082031 -6.363281 C 3.816406 -6.363281 4.421875 -6.066406 4.898438 -5.472656 L 4.898438 -6.222656 L 5.871094 -6.222656 L 5.871094 -0.84375 C 5.871094 0.125 5.769531 0.808594 5.574219 1.214844 C 5.375 1.613281 5.0625 1.933594 4.636719 2.171875 C 4.207031 2.402344 3.683594 2.519531 3.058594 2.523438 C 2.316406 2.519531 1.714844 2.351563 1.257813 2.023438 C 0.800781 1.6875 0.582031 1.1875 0.597656 0.515625 Z M 1.46875 -3.222656 C 1.464844 -2.40625 1.628906 -1.808594 1.957031 -1.4375 C 2.28125 -1.058594 2.6875 -0.871094 3.175781 -0.875 C 3.660156 -0.871094 4.066406 -1.058594 4.394531 -1.433594 C 4.722656 -1.804688 4.886719 -2.390625 4.886719 -3.1875 C 4.886719 -3.945313 4.714844 -4.519531 4.378906 -4.910156 C 4.039063 -5.296875 3.632813 -5.488281 3.15625 -5.492188 C 2.683594 -5.488281 2.285156 -5.296875 1.960938 -4.917969 C 1.628906 -4.535156 1.464844 -3.972656 1.46875 -3.222656 Z M 1.46875 -3.222656 "/>
</symbol>
<symbol overflow="visible" id="glyph1-7">
<path style="stroke:none;" d="M -0.179688 2.382813 L -0.179688 1.625 L 6.808594 1.625 L 6.808594 2.382813 Z M -0.179688 2.382813 "/>
</symbol>
<symbol overflow="visible" id="glyph1-8">
<path style="stroke:none;" d="M 0.914063 0 L 0.914063 -8.589844 L 2.078125 -8.589844 L 6.59375 -1.84375 L 6.59375 -8.589844 L 7.679688 -8.589844 L 7.679688 0 L 6.515625 0 L 2.003906 -6.75 L 2.003906 0 Z M 0.914063 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-9">
<path style="stroke:none;" d="M 4.867188 0 L 4.867188 -0.914063 C 4.378906 -0.210938 3.722656 0.140625 2.894531 0.140625 C 2.527344 0.140625 2.183594 0.0703125 1.867188 -0.0703125 C 1.546875 -0.210938 1.308594 -0.386719 1.15625 -0.601563 C 1 -0.8125 0.894531 -1.074219 0.832031 -1.382813 C 0.785156 -1.589844 0.761719 -1.917969 0.765625 -2.367188 L 0.765625 -6.222656 L 1.820313 -6.222656 L 1.820313 -2.773438 C 1.816406 -2.21875 1.839844 -1.847656 1.886719 -1.65625 C 1.949219 -1.378906 2.089844 -1.160156 2.308594 -1.003906 C 2.523438 -0.839844 2.789063 -0.761719 3.105469 -0.765625 C 3.417969 -0.761719 3.714844 -0.84375 3.996094 -1.007813 C 4.273438 -1.171875 4.46875 -1.390625 4.585938 -1.671875 C 4.699219 -1.949219 4.757813 -2.355469 4.757813 -2.890625 L 4.757813 -6.222656 L 5.8125 -6.222656 L 5.8125 0 Z M 4.867188 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-10">
<path style="stroke:none;" d="M 0.789063 0 L 0.789063 -6.222656 L 1.734375 -6.222656 L 1.734375 -5.351563 C 1.929688 -5.648438 2.1875 -5.894531 2.511719 -6.082031 C 2.835938 -6.269531 3.207031 -6.363281 3.621094 -6.363281 C 4.082031 -6.363281 4.457031 -6.265625 4.753906 -6.074219 C 5.042969 -5.882813 5.253906 -5.617188 5.378906 -5.273438 C 5.871094 -6 6.511719 -6.363281 7.300781 -6.363281 C 7.917969 -6.363281 8.390625 -6.191406 8.722656 -5.847656 C 9.054688 -5.503906 9.222656 -4.976563 9.222656 -4.273438 L 9.222656 0 L 8.171875 0 L 8.171875 -3.921875 C 8.167969 -4.339844 8.132813 -4.644531 8.070313 -4.832031 C 8 -5.015625 7.878906 -5.164063 7.699219 -5.277344 C 7.519531 -5.390625 7.308594 -5.449219 7.066406 -5.449219 C 6.628906 -5.449219 6.265625 -5.300781 5.976563 -5.011719 C 5.6875 -4.71875 5.542969 -4.253906 5.542969 -3.617188 L 5.542969 0 L 4.488281 0 L 4.488281 -4.042969 C 4.488281 -4.511719 4.402344 -4.863281 4.230469 -5.097656 C 4.058594 -5.332031 3.777344 -5.449219 3.386719 -5.449219 C 3.089844 -5.449219 2.8125 -5.371094 2.5625 -5.214844 C 2.308594 -5.058594 2.128906 -4.828125 2.015625 -4.527344 C 1.898438 -4.226563 1.839844 -3.792969 1.84375 -3.226563 L 1.84375 0 Z M 0.789063 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-11">
<path style="stroke:none;" d="M 1.765625 0 L 0.785156 0 L 0.785156 -8.589844 L 1.839844 -8.589844 L 1.839844 -5.523438 C 2.285156 -6.082031 2.851563 -6.363281 3.546875 -6.363281 C 3.921875 -6.363281 4.285156 -6.285156 4.628906 -6.128906 C 4.972656 -5.972656 5.253906 -5.753906 5.472656 -5.480469 C 5.691406 -5.199219 5.863281 -4.863281 5.992188 -4.46875 C 6.113281 -4.074219 6.175781 -3.652344 6.179688 -3.203125 C 6.175781 -2.136719 5.914063 -1.3125 5.390625 -0.730469 C 4.863281 -0.148438 4.230469 0.140625 3.492188 0.140625 C 2.757813 0.140625 2.179688 -0.164063 1.765625 -0.78125 Z M 1.75 -3.15625 C 1.746094 -2.410156 1.847656 -1.871094 2.054688 -1.539063 C 2.386719 -0.996094 2.835938 -0.726563 3.40625 -0.726563 C 3.859375 -0.726563 4.257813 -0.925781 4.597656 -1.328125 C 4.929688 -1.726563 5.097656 -2.324219 5.101563 -3.117188 C 5.097656 -3.929688 4.9375 -4.527344 4.617188 -4.914063 C 4.296875 -5.300781 3.90625 -5.496094 3.453125 -5.496094 C 2.984375 -5.496094 2.585938 -5.292969 2.253906 -4.894531 C 1.914063 -4.492188 1.746094 -3.914063 1.75 -3.15625 Z M 1.75 -3.15625 "/>
</symbol>
<symbol overflow="visible" id="glyph1-12">
<path style="stroke:none;" d="M 0.578125 -4.183594 C 0.574219 -5.605469 0.957031 -6.71875 1.726563 -7.53125 C 2.488281 -8.335938 3.476563 -8.742188 4.695313 -8.742188 C 5.484375 -8.742188 6.199219 -8.550781 6.835938 -8.171875 C 7.472656 -7.792969 7.957031 -7.265625 8.292969 -6.585938 C 8.625 -5.90625 8.792969 -5.136719 8.796875 -4.28125 C 8.792969 -3.410156 8.617188 -2.632813 8.269531 -1.945313 C 7.914063 -1.257813 7.417969 -0.734375 6.773438 -0.382813 C 6.125 -0.0273438 5.429688 0.144531 4.6875 0.148438 C 3.878906 0.144531 3.15625 -0.046875 2.519531 -0.4375 C 1.878906 -0.824219 1.394531 -1.359375 1.070313 -2.039063 C 0.738281 -2.714844 0.574219 -3.429688 0.578125 -4.183594 Z M 1.75 -4.164063 C 1.746094 -3.128906 2.023438 -2.3125 2.585938 -1.71875 C 3.140625 -1.121094 3.839844 -0.824219 4.679688 -0.828125 C 5.535156 -0.824219 6.238281 -1.125 6.792969 -1.730469 C 7.34375 -2.328125 7.621094 -3.183594 7.625 -4.289063 C 7.621094 -4.984375 7.503906 -5.59375 7.269531 -6.117188 C 7.03125 -6.640625 6.683594 -7.042969 6.230469 -7.332031 C 5.769531 -7.617188 5.261719 -7.761719 4.699219 -7.765625 C 3.894531 -7.761719 3.199219 -7.484375 2.621094 -6.933594 C 2.035156 -6.378906 1.746094 -5.457031 1.75 -4.164063 Z M 1.75 -4.164063 "/>
</symbol>
<symbol overflow="visible" id="glyph1-13">
<path style="stroke:none;" d="M 1.042969 0 L 1.042969 -5.402344 L 0.109375 -5.402344 L 0.109375 -6.222656 L 1.042969 -6.222656 L 1.042969 -6.882813 C 1.042969 -7.300781 1.078125 -7.613281 1.15625 -7.816406 C 1.25 -8.089844 1.429688 -8.308594 1.6875 -8.480469 C 1.945313 -8.644531 2.304688 -8.730469 2.765625 -8.734375 C 3.0625 -8.730469 3.390625 -8.695313 3.75 -8.632813 L 3.59375 -7.710938 C 3.371094 -7.75 3.164063 -7.769531 2.96875 -7.769531 C 2.648438 -7.769531 2.421875 -7.699219 2.292969 -7.5625 C 2.15625 -7.425781 2.089844 -7.171875 2.09375 -6.796875 L 2.09375 -6.222656 L 3.304688 -6.222656 L 3.304688 -5.402344 L 2.09375 -5.402344 L 2.09375 0 Z M 1.042969 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-14">
<path style="stroke:none;" d="M 7.054688 -3.011719 L 8.191406 -2.726563 C 7.953125 -1.789063 7.523438 -1.078125 6.90625 -0.585938 C 6.285156 -0.0976563 5.527344 0.144531 4.632813 0.148438 C 3.707031 0.144531 2.953125 -0.0390625 2.375 -0.417969 C 1.792969 -0.792969 1.351563 -1.339844 1.050781 -2.054688 C 0.746094 -2.769531 0.597656 -3.539063 0.597656 -4.359375 C 0.597656 -5.253906 0.765625 -6.03125 1.109375 -6.699219 C 1.449219 -7.363281 1.9375 -7.871094 2.570313 -8.214844 C 3.199219 -8.558594 3.894531 -8.730469 4.652344 -8.734375 C 5.511719 -8.730469 6.234375 -8.511719 6.820313 -8.078125 C 7.40625 -7.636719 7.8125 -7.023438 8.046875 -6.234375 L 6.925781 -5.96875 C 6.722656 -6.589844 6.433594 -7.046875 6.058594 -7.335938 C 5.679688 -7.621094 5.203125 -7.761719 4.628906 -7.765625 C 3.96875 -7.761719 3.414063 -7.605469 2.972656 -7.289063 C 2.527344 -6.96875 2.21875 -6.542969 2.039063 -6.011719 C 1.859375 -5.480469 1.769531 -4.929688 1.769531 -4.367188 C 1.769531 -3.632813 1.875 -2.996094 2.085938 -2.449219 C 2.296875 -1.902344 2.628906 -1.496094 3.082031 -1.230469 C 3.53125 -0.960938 4.015625 -0.824219 4.539063 -0.828125 C 5.175781 -0.824219 5.714844 -1.007813 6.15625 -1.378906 C 6.597656 -1.742188 6.898438 -2.289063 7.054688 -3.011719 Z M 7.054688 -3.011719 "/>
</symbol>
<symbol overflow="visible" id="glyph1-15">
<path style="stroke:none;" d="M 0.789063 0 L 0.789063 -8.589844 L 1.84375 -8.589844 L 1.84375 -5.507813 C 2.335938 -6.078125 2.957031 -6.363281 3.710938 -6.363281 C 4.164063 -6.363281 4.566406 -6.269531 4.910156 -6.089844 C 5.25 -5.90625 5.492188 -5.65625 5.640625 -5.339844 C 5.785156 -5.015625 5.859375 -4.550781 5.859375 -3.945313 L 5.859375 0 L 4.804688 0 L 4.804688 -3.945313 C 4.804688 -4.46875 4.6875 -4.851563 4.460938 -5.09375 C 4.226563 -5.328125 3.90625 -5.449219 3.492188 -5.453125 C 3.179688 -5.449219 2.882813 -5.367188 2.609375 -5.210938 C 2.328125 -5.046875 2.132813 -4.828125 2.019531 -4.550781 C 1.898438 -4.273438 1.839844 -3.890625 1.84375 -3.40625 L 1.84375 0 Z M 0.789063 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-16">
<path style="stroke:none;" d="M 0.796875 -7.375 L 0.796875 -8.589844 L 1.851563 -8.589844 L 1.851563 -7.375 Z M 0.796875 0 L 0.796875 -6.222656 L 1.851563 -6.222656 L 1.851563 0 Z M 0.796875 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-17">
<path style="stroke:none;" d="M 0.765625 0 L 0.765625 -8.589844 L 1.820313 -8.589844 L 1.820313 0 Z M 0.765625 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-18">
<path style="stroke:none;" d="M 4.828125 0 L 4.828125 -0.785156 C 4.429688 -0.167969 3.847656 0.140625 3.085938 0.140625 C 2.589844 0.140625 2.132813 0.00390625 1.71875 -0.269531 C 1.296875 -0.542969 0.976563 -0.921875 0.75 -1.414063 C 0.523438 -1.898438 0.410156 -2.464844 0.410156 -3.105469 C 0.410156 -3.726563 0.511719 -4.289063 0.71875 -4.796875 C 0.925781 -5.300781 1.238281 -5.6875 1.652344 -5.957031 C 2.066406 -6.226563 2.527344 -6.363281 3.039063 -6.363281 C 3.410156 -6.363281 3.746094 -6.28125 4.042969 -6.125 C 4.335938 -5.964844 4.574219 -5.761719 4.757813 -5.507813 L 4.757813 -8.589844 L 5.804688 -8.589844 L 5.804688 0 Z M 1.492188 -3.105469 C 1.488281 -2.308594 1.65625 -1.710938 1.996094 -1.316406 C 2.328125 -0.921875 2.726563 -0.726563 3.1875 -0.726563 C 3.648438 -0.726563 4.039063 -0.914063 4.359375 -1.292969 C 4.679688 -1.667969 4.839844 -2.242188 4.84375 -3.015625 C 4.839844 -3.867188 4.675781 -4.492188 4.351563 -4.894531 C 4.019531 -5.289063 3.617188 -5.488281 3.140625 -5.492188 C 2.671875 -5.488281 2.277344 -5.296875 1.964844 -4.917969 C 1.644531 -4.53125 1.488281 -3.929688 1.492188 -3.105469 Z M 1.492188 -3.105469 "/>
</symbol>
<symbol overflow="visible" id="glyph1-19">
<path style="stroke:none;" d="M 0.789063 0 L 0.789063 -6.222656 L 1.742188 -6.222656 L 1.742188 -5.335938 C 2.195313 -6.019531 2.855469 -6.363281 3.71875 -6.363281 C 4.089844 -6.363281 4.433594 -6.292969 4.753906 -6.160156 C 5.066406 -6.023438 5.304688 -5.847656 5.460938 -5.632813 C 5.617188 -5.410156 5.726563 -5.152344 5.789063 -4.851563 C 5.828125 -4.65625 5.847656 -4.3125 5.847656 -3.828125 L 5.847656 0 L 4.792969 0 L 4.792969 -3.785156 C 4.792969 -4.214844 4.75 -4.535156 4.667969 -4.75 C 4.585938 -4.960938 4.441406 -5.128906 4.234375 -5.257813 C 4.023438 -5.382813 3.777344 -5.449219 3.5 -5.449219 C 3.046875 -5.449219 2.660156 -5.304688 2.332031 -5.019531 C 2.003906 -4.734375 1.839844 -4.195313 1.84375 -3.398438 L 1.84375 0 Z M 0.789063 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-20">
<path style="stroke:none;" d="M 0.925781 0 L 0.925781 -8.589844 L 4.164063 -8.589844 C 4.734375 -8.589844 5.171875 -8.5625 5.472656 -8.507813 C 5.894531 -8.4375 6.246094 -8.300781 6.53125 -8.105469 C 6.816406 -7.90625 7.046875 -7.632813 7.222656 -7.277344 C 7.394531 -6.917969 7.480469 -6.527344 7.484375 -6.105469 C 7.480469 -5.371094 7.25 -4.75 6.785156 -4.25 C 6.316406 -3.742188 5.476563 -3.492188 4.265625 -3.492188 L 2.0625 -3.492188 L 2.0625 0 Z M 2.0625 -4.507813 L 4.28125 -4.507813 C 5.011719 -4.503906 5.535156 -4.640625 5.847656 -4.917969 C 6.15625 -5.1875 6.308594 -5.574219 6.3125 -6.070313 C 6.308594 -6.429688 6.21875 -6.734375 6.039063 -6.992188 C 5.855469 -7.242188 5.617188 -7.414063 5.320313 -7.5 C 5.125 -7.550781 4.769531 -7.574219 4.257813 -7.578125 L 2.0625 -7.578125 Z M 2.0625 -4.507813 "/>
</symbol>
<symbol overflow="visible" id="glyph1-21">
<path style="stroke:none;" d="M 0.878906 0 L 0.878906 -8.589844 L 4.101563 -8.589844 C 4.757813 -8.589844 5.28125 -8.5 5.679688 -8.328125 C 6.070313 -8.152344 6.382813 -7.886719 6.609375 -7.527344 C 6.835938 -7.164063 6.949219 -6.785156 6.949219 -6.390625 C 6.949219 -6.023438 6.847656 -5.679688 6.648438 -5.355469 C 6.449219 -5.027344 6.148438 -4.765625 5.75 -4.570313 C 6.265625 -4.417969 6.664063 -4.15625 6.945313 -3.792969 C 7.222656 -3.421875 7.363281 -2.988281 7.367188 -2.492188 C 7.363281 -2.085938 7.277344 -1.710938 7.109375 -1.367188 C 6.9375 -1.019531 6.730469 -0.753906 6.480469 -0.570313 C 6.230469 -0.378906 5.914063 -0.238281 5.539063 -0.144531 C 5.160156 -0.046875 4.699219 0 4.15625 0 Z M 2.015625 -4.980469 L 3.875 -4.980469 C 4.375 -4.980469 4.738281 -5.011719 4.957031 -5.078125 C 5.246094 -5.164063 5.460938 -5.308594 5.609375 -5.507813 C 5.75 -5.703125 5.824219 -5.953125 5.828125 -6.257813 C 5.824219 -6.542969 5.757813 -6.792969 5.625 -7.011719 C 5.488281 -7.226563 5.292969 -7.375 5.039063 -7.457031 C 4.78125 -7.535156 4.34375 -7.574219 3.734375 -7.578125 L 2.015625 -7.578125 Z M 2.015625 -1.015625 L 4.15625 -1.015625 C 4.515625 -1.011719 4.773438 -1.027344 4.929688 -1.054688 C 5.1875 -1.101563 5.40625 -1.179688 5.582031 -1.289063 C 5.757813 -1.398438 5.902344 -1.554688 6.015625 -1.765625 C 6.128906 -1.96875 6.1875 -2.210938 6.1875 -2.492188 C 6.1875 -2.804688 6.105469 -3.082031 5.941406 -3.324219 C 5.777344 -3.558594 5.546875 -3.726563 5.257813 -3.824219 C 4.960938 -3.917969 4.542969 -3.964844 4 -3.96875 L 2.015625 -3.96875 Z M 2.015625 -1.015625 "/>
</symbol>
<symbol overflow="visible" id="glyph1-22">
<path style="stroke:none;" d="M 0.367188 -1.859375 L 1.414063 -2.023438 C 1.46875 -1.601563 1.632813 -1.28125 1.902344 -1.058594 C 2.167969 -0.835938 2.542969 -0.726563 3.023438 -0.726563 C 3.507813 -0.726563 3.867188 -0.824219 4.101563 -1.023438 C 4.335938 -1.21875 4.453125 -1.449219 4.453125 -1.71875 C 4.453125 -1.953125 4.347656 -2.140625 4.140625 -2.28125 C 3.996094 -2.371094 3.636719 -2.492188 3.0625 -2.636719 C 2.289063 -2.832031 1.753906 -3 1.457031 -3.144531 C 1.15625 -3.285156 0.929688 -3.480469 0.777344 -3.734375 C 0.621094 -3.984375 0.542969 -4.265625 0.546875 -4.570313 C 0.542969 -4.84375 0.605469 -5.097656 0.734375 -5.339844 C 0.859375 -5.574219 1.035156 -5.773438 1.253906 -5.929688 C 1.417969 -6.046875 1.640625 -6.148438 1.925781 -6.234375 C 2.207031 -6.320313 2.511719 -6.363281 2.835938 -6.363281 C 3.324219 -6.363281 3.75 -6.292969 4.121094 -6.152344 C 4.488281 -6.011719 4.761719 -5.820313 4.9375 -5.578125 C 5.113281 -5.335938 5.234375 -5.015625 5.304688 -4.617188 L 4.273438 -4.476563 C 4.222656 -4.796875 4.085938 -5.046875 3.863281 -5.226563 C 3.636719 -5.40625 3.320313 -5.496094 2.914063 -5.496094 C 2.425781 -5.496094 2.082031 -5.414063 1.875 -5.253906 C 1.664063 -5.09375 1.558594 -4.90625 1.5625 -4.695313 C 1.558594 -4.554688 1.601563 -4.433594 1.695313 -4.324219 C 1.773438 -4.210938 1.910156 -4.117188 2.097656 -4.042969 C 2.203125 -4.003906 2.511719 -3.914063 3.03125 -3.773438 C 3.773438 -3.574219 4.292969 -3.410156 4.589844 -3.285156 C 4.878906 -3.15625 5.113281 -2.972656 5.285156 -2.730469 C 5.453125 -2.488281 5.535156 -2.1875 5.539063 -1.828125 C 5.535156 -1.476563 5.433594 -1.144531 5.230469 -0.832031 C 5.023438 -0.519531 4.726563 -0.277344 4.339844 -0.113281 C 3.953125 0.0585938 3.515625 0.140625 3.03125 0.140625 C 2.21875 0.140625 1.601563 -0.0273438 1.179688 -0.363281 C 0.753906 -0.699219 0.484375 -1.195313 0.367188 -1.859375 Z M 0.367188 -1.859375 "/>
</symbol>
<symbol overflow="visible" id="glyph1-23">
<path style="stroke:none;" d="M 0.5 -4.234375 C 0.496094 -5.246094 0.601563 -6.0625 0.8125 -6.6875 C 1.019531 -7.304688 1.328125 -7.785156 1.742188 -8.121094 C 2.148438 -8.457031 2.667969 -8.625 3.296875 -8.625 C 3.757813 -8.625 4.164063 -8.53125 4.511719 -8.347656 C 4.855469 -8.160156 5.140625 -7.890625 5.371094 -7.542969 C 5.59375 -7.191406 5.773438 -6.765625 5.90625 -6.265625 C 6.035156 -5.761719 6.097656 -5.085938 6.101563 -4.234375 C 6.097656 -3.226563 5.996094 -2.414063 5.789063 -1.796875 C 5.578125 -1.175781 5.265625 -0.695313 4.859375 -0.359375 C 4.445313 -0.0195313 3.925781 0.144531 3.296875 0.148438 C 2.464844 0.144531 1.816406 -0.148438 1.347656 -0.742188 C 0.78125 -1.457031 0.496094 -2.621094 0.5 -4.234375 Z M 1.582031 -4.234375 C 1.582031 -2.824219 1.746094 -1.886719 2.074219 -1.417969 C 2.402344 -0.949219 2.808594 -0.714844 3.296875 -0.71875 C 3.777344 -0.714844 4.183594 -0.949219 4.519531 -1.421875 C 4.847656 -1.886719 5.015625 -2.824219 5.015625 -4.234375 C 5.015625 -5.648438 4.847656 -6.589844 4.519531 -7.054688 C 4.183594 -7.515625 3.773438 -7.746094 3.289063 -7.75 C 2.800781 -7.746094 2.414063 -7.542969 2.125 -7.136719 C 1.761719 -6.613281 1.582031 -5.644531 1.582031 -4.234375 Z M 1.582031 -4.234375 "/>
</symbol>
<symbol overflow="visible" id="glyph1-24">
<path style="stroke:none;" d="M 1.089844 0 L 1.089844 -1.203125 L 2.289063 -1.203125 L 2.289063 0 Z M 1.089844 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-25">
<path style="stroke:none;" d="M 0.5 -2.25 L 1.605469 -2.34375 C 1.683594 -1.804688 1.871094 -1.398438 2.175781 -1.125 C 2.472656 -0.851563 2.835938 -0.714844 3.257813 -0.71875 C 3.765625 -0.714844 4.195313 -0.90625 4.546875 -1.292969 C 4.898438 -1.671875 5.074219 -2.179688 5.074219 -2.820313 C 5.074219 -3.414063 4.902344 -3.890625 4.566406 -4.242188 C 4.226563 -4.589844 3.785156 -4.761719 3.242188 -4.765625 C 2.898438 -4.761719 2.59375 -4.683594 2.320313 -4.53125 C 2.046875 -4.375 1.832031 -4.175781 1.675781 -3.929688 L 0.6875 -4.0625 L 1.515625 -8.472656 L 5.789063 -8.472656 L 5.789063 -7.464844 L 2.359375 -7.464844 L 1.898438 -5.15625 C 2.414063 -5.515625 2.953125 -5.695313 3.523438 -5.695313 C 4.269531 -5.695313 4.902344 -5.433594 5.421875 -4.914063 C 5.933594 -4.394531 6.191406 -3.726563 6.195313 -2.914063 C 6.191406 -2.132813 5.964844 -1.460938 5.515625 -0.898438 C 4.960938 -0.199219 4.210938 0.144531 3.257813 0.148438 C 2.476563 0.144531 1.835938 -0.0703125 1.34375 -0.507813 C 0.84375 -0.941406 0.5625 -1.523438 0.5 -2.25 Z M 0.5 -2.25 "/>
</symbol>
<symbol overflow="visible" id="glyph1-26">
<path style="stroke:none;" d="M 5.96875 -6.484375 L 4.921875 -6.40625 C 4.828125 -6.8125 4.695313 -7.113281 4.523438 -7.304688 C 4.234375 -7.605469 3.882813 -7.757813 3.46875 -7.757813 C 3.132813 -7.757813 2.835938 -7.664063 2.585938 -7.476563 C 2.25 -7.234375 1.988281 -6.878906 1.796875 -6.414063 C 1.605469 -5.949219 1.507813 -5.289063 1.5 -4.429688 C 1.753906 -4.8125 2.0625 -5.097656 2.433594 -5.289063 C 2.796875 -5.472656 3.183594 -5.566406 3.585938 -5.570313 C 4.289063 -5.566406 4.886719 -5.308594 5.382813 -4.792969 C 5.875 -4.277344 6.121094 -3.609375 6.125 -2.789063 C 6.121094 -2.25 6.003906 -1.746094 5.773438 -1.285156 C 5.539063 -0.820313 5.222656 -0.46875 4.816406 -0.222656 C 4.410156 0.0234375 3.949219 0.144531 3.433594 0.148438 C 2.554688 0.144531 1.835938 -0.175781 1.285156 -0.820313 C 0.726563 -1.46875 0.449219 -2.535156 0.453125 -4.019531 C 0.449219 -5.675781 0.757813 -6.882813 1.371094 -7.640625 C 1.902344 -8.296875 2.621094 -8.625 3.53125 -8.625 C 4.207031 -8.625 4.761719 -8.433594 5.195313 -8.054688 C 5.625 -7.675781 5.882813 -7.152344 5.96875 -6.484375 Z M 1.664063 -2.78125 C 1.664063 -2.417969 1.738281 -2.070313 1.894531 -1.738281 C 2.042969 -1.40625 2.261719 -1.152344 2.542969 -0.980469 C 2.820313 -0.800781 3.109375 -0.714844 3.414063 -0.71875 C 3.859375 -0.714844 4.242188 -0.894531 4.566406 -1.257813 C 4.882813 -1.613281 5.042969 -2.101563 5.046875 -2.726563 C 5.042969 -3.316406 4.886719 -3.785156 4.570313 -4.128906 C 4.25 -4.46875 3.851563 -4.640625 3.375 -4.640625 C 2.898438 -4.640625 2.492188 -4.46875 2.160156 -4.128906 C 1.828125 -3.785156 1.664063 -3.335938 1.664063 -2.78125 Z M 1.664063 -2.78125 "/>
</symbol>
<symbol overflow="visible" id="glyph1-27">
<path style="stroke:none;" d="M 0.570313 -7.464844 L 0.570313 -8.476563 L 6.128906 -8.476563 L 6.128906 -7.65625 C 5.582031 -7.074219 5.039063 -6.300781 4.5 -5.335938 C 3.960938 -4.371094 3.546875 -3.378906 3.257813 -2.359375 C 3.046875 -1.636719 2.910156 -0.851563 2.851563 0 L 1.769531 0 C 1.78125 -0.675781 1.914063 -1.492188 2.167969 -2.449219 C 2.417969 -3.402344 2.78125 -4.324219 3.257813 -5.214844 C 3.734375 -6.105469 4.238281 -6.855469 4.773438 -7.464844 Z M 0.570313 -7.464844 "/>
</symbol>
<symbol overflow="visible" id="glyph1-28">
<path style="stroke:none;" d="M 2.121094 -4.65625 C 1.683594 -4.816406 1.359375 -5.046875 1.148438 -5.34375 C 0.9375 -5.640625 0.832031 -5.996094 0.832031 -6.410156 C 0.832031 -7.035156 1.054688 -7.558594 1.503906 -7.984375 C 1.953125 -8.410156 2.550781 -8.625 3.296875 -8.625 C 4.042969 -8.625 4.648438 -8.40625 5.109375 -7.972656 C 5.566406 -7.535156 5.792969 -7.003906 5.796875 -6.382813 C 5.792969 -5.976563 5.6875 -5.628906 5.480469 -5.339844 C 5.269531 -5.042969 4.953125 -4.816406 4.53125 -4.65625 C 5.054688 -4.480469 5.457031 -4.203125 5.734375 -3.824219 C 6.007813 -3.4375 6.144531 -2.980469 6.148438 -2.453125 C 6.144531 -1.714844 5.886719 -1.097656 5.367188 -0.601563 C 4.84375 -0.101563 4.160156 0.144531 3.316406 0.148438 C 2.46875 0.144531 1.785156 -0.101563 1.265625 -0.605469 C 0.742188 -1.105469 0.480469 -1.734375 0.484375 -2.484375 C 0.480469 -3.039063 0.621094 -3.503906 0.910156 -3.886719 C 1.191406 -4.261719 1.597656 -4.519531 2.121094 -4.65625 Z M 1.910156 -6.445313 C 1.910156 -6.039063 2.039063 -5.707031 2.300781 -5.449219 C 2.5625 -5.191406 2.902344 -5.0625 3.320313 -5.0625 C 3.722656 -5.0625 4.054688 -5.1875 4.320313 -5.445313 C 4.578125 -5.695313 4.710938 -6.011719 4.710938 -6.386719 C 4.710938 -6.773438 4.574219 -7.097656 4.308594 -7.363281 C 4.035156 -7.625 3.703125 -7.757813 3.3125 -7.757813 C 2.90625 -7.757813 2.574219 -7.628906 2.308594 -7.371094 C 2.042969 -7.113281 1.910156 -6.804688 1.910156 -6.445313 Z M 1.570313 -2.476563 C 1.570313 -2.175781 1.640625 -1.886719 1.785156 -1.605469 C 1.925781 -1.324219 2.136719 -1.105469 2.421875 -0.949219 C 2.699219 -0.792969 3.003906 -0.714844 3.328125 -0.71875 C 3.832031 -0.714844 4.246094 -0.878906 4.578125 -1.207031 C 4.902344 -1.53125 5.066406 -1.941406 5.070313 -2.445313 C 5.066406 -2.945313 4.898438 -3.367188 4.5625 -3.703125 C 4.222656 -4.035156 3.800781 -4.199219 3.292969 -4.203125 C 2.792969 -4.199219 2.378906 -4.035156 2.058594 -3.710938 C 1.730469 -3.378906 1.570313 -2.96875 1.570313 -2.476563 Z M 1.570313 -2.476563 "/>
</symbol>
<symbol overflow="visible" id="glyph1-29">
<path style="stroke:none;" d="M 0.65625 -1.984375 L 1.671875 -2.078125 C 1.75 -1.601563 1.914063 -1.257813 2.160156 -1.042969 C 2.398438 -0.824219 2.710938 -0.714844 3.09375 -0.71875 C 3.414063 -0.714844 3.695313 -0.789063 3.945313 -0.941406 C 4.1875 -1.085938 4.390625 -1.285156 4.546875 -1.535156 C 4.703125 -1.785156 4.832031 -2.121094 4.9375 -2.542969 C 5.042969 -2.964844 5.097656 -3.394531 5.097656 -3.832031 C 5.097656 -3.878906 5.09375 -3.949219 5.09375 -4.042969 C 4.875 -3.707031 4.585938 -3.433594 4.226563 -3.226563 C 3.859375 -3.015625 3.464844 -2.910156 3.039063 -2.914063 C 2.328125 -2.910156 1.726563 -3.167969 1.238281 -3.6875 C 0.742188 -4.199219 0.496094 -4.878906 0.5 -5.726563 C 0.496094 -6.59375 0.753906 -7.296875 1.269531 -7.828125 C 1.78125 -8.359375 2.425781 -8.625 3.199219 -8.625 C 3.757813 -8.625 4.265625 -8.472656 4.730469 -8.171875 C 5.191406 -7.871094 5.542969 -7.441406 5.785156 -6.886719 C 6.023438 -6.328125 6.144531 -5.523438 6.148438 -4.46875 C 6.144531 -3.371094 6.027344 -2.496094 5.789063 -1.847656 C 5.546875 -1.195313 5.191406 -0.703125 4.722656 -0.363281 C 4.253906 -0.0234375 3.703125 0.144531 3.070313 0.148438 C 2.398438 0.144531 1.847656 -0.0390625 1.421875 -0.410156 C 0.996094 -0.785156 0.742188 -1.308594 0.65625 -1.984375 Z M 4.976563 -5.777344 C 4.972656 -6.382813 4.8125 -6.863281 4.492188 -7.21875 C 4.167969 -7.570313 3.78125 -7.746094 3.328125 -7.75 C 2.859375 -7.746094 2.449219 -7.554688 2.101563 -7.175781 C 1.753906 -6.789063 1.582031 -6.292969 1.582031 -5.6875 C 1.582031 -5.136719 1.746094 -4.691406 2.074219 -4.355469 C 2.402344 -4.011719 2.808594 -3.84375 3.296875 -3.84375 C 3.785156 -3.84375 4.1875 -4.011719 4.503906 -4.355469 C 4.816406 -4.691406 4.972656 -5.167969 4.976563 -5.777344 Z M 4.976563 -5.777344 "/>
</symbol>
<symbol overflow="visible" id="glyph1-30">
<path style="stroke:none;" d="M 4.46875 0 L 3.414063 0 L 3.414063 -6.71875 C 3.160156 -6.476563 2.828125 -6.234375 2.414063 -5.996094 C 2 -5.75 1.628906 -5.570313 1.304688 -5.449219 L 1.304688 -6.46875 C 1.894531 -6.742188 2.410156 -7.078125 2.851563 -7.476563 C 3.292969 -7.871094 3.605469 -8.253906 3.789063 -8.625 L 4.46875 -8.625 Z M 4.46875 0 "/>
</symbol>
<symbol overflow="visible" id="glyph2-0">
<path style="stroke:none;" d="M 0 -1.5 L -7.5 -1.5 L -7.5 -7.5 L 0 -7.5 Z M -0.1875 -1.6875 L -0.1875 -7.3125 L -7.3125 -7.3125 L -7.3125 -1.6875 Z M -0.1875 -1.6875 "/>
</symbol>
<symbol overflow="visible" id="glyph2-1">
<path style="stroke:none;" d="M 0 -0.984375 L -8.589844 -0.984375 L -8.589844 -6.78125 L -7.578125 -6.78125 L -7.578125 -2.121094 L -4.914063 -2.121094 L -4.914063 -6.152344 L -3.902344 -6.152344 L -3.902344 -2.121094 L 0 -2.121094 Z M 0 -0.984375 "/>
</symbol>
<symbol overflow="visible" id="glyph2-2">
<path style="stroke:none;" d="M 0 -0.78125 L -6.222656 -0.78125 L -6.222656 -1.730469 L -5.28125 -1.730469 C -5.71875 -1.96875 -6.011719 -2.191406 -6.152344 -2.398438 C -6.292969 -2.601563 -6.363281 -2.828125 -6.363281 -3.078125 C -6.363281 -3.429688 -6.25 -3.792969 -6.023438 -4.160156 L -5.046875 -3.796875 C -5.195313 -3.539063 -5.273438 -3.28125 -5.273438 -3.023438 C -5.273438 -2.792969 -5.203125 -2.585938 -5.066406 -2.402344 C -4.925781 -2.21875 -4.734375 -2.085938 -4.488281 -2.011719 C -4.113281 -1.890625 -3.703125 -1.832031 -3.257813 -1.835938 L 0 -1.835938 Z M 0 -0.78125 "/>
</symbol>
<symbol overflow="visible" id="glyph2-3">
<path style="stroke:none;" d="M -2.003906 -5.050781 L -1.867188 -6.140625 C -1.230469 -5.96875 -0.738281 -5.648438 -0.386719 -5.183594 C -0.0351563 -4.71875 0.140625 -4.125 0.140625 -3.40625 C 0.140625 -2.492188 -0.136719 -1.769531 -0.699219 -1.238281 C -1.253906 -0.703125 -2.042969 -0.4375 -3.058594 -0.441406 C -4.105469 -0.4375 -4.917969 -0.707031 -5.496094 -1.25 C -6.074219 -1.785156 -6.363281 -2.484375 -6.363281 -3.347656 C -6.363281 -4.175781 -6.078125 -4.855469 -5.511719 -5.382813 C -4.945313 -5.910156 -4.148438 -6.175781 -3.121094 -6.175781 C -3.054688 -6.175781 -2.960938 -6.171875 -2.839844 -6.171875 L -2.84375 -1.53125 C -2.15625 -1.566406 -1.632813 -1.761719 -1.269531 -2.109375 C -0.90625 -2.457031 -0.726563 -2.890625 -0.726563 -3.410156 C -0.726563 -3.796875 -0.828125 -4.125 -1.03125 -4.402344 C -1.234375 -4.671875 -1.558594 -4.890625 -2.003906 -5.050781 Z M -3.710938 -1.589844 L -3.707031 -5.0625 C -4.226563 -5.015625 -4.621094 -4.882813 -4.886719 -4.664063 C -5.292969 -4.328125 -5.496094 -3.890625 -5.496094 -3.359375 C -5.496094 -2.871094 -5.332031 -2.464844 -5.007813 -2.136719 C -4.683594 -1.804688 -4.25 -1.621094 -3.710938 -1.589844 Z M -3.710938 -1.589844 "/>
</symbol>
<symbol overflow="visible" id="glyph2-4">
<path style="stroke:none;" d="M 2.386719 -4.757813 L -0.660156 -4.757813 C -0.429688 -4.59375 -0.238281 -4.363281 -0.0859375 -4.066406 C 0.0664063 -3.769531 0.140625 -3.457031 0.140625 -3.128906 C 0.140625 -2.390625 -0.152344 -1.753906 -0.742188 -1.222656 C -1.332031 -0.6875 -2.140625 -0.421875 -3.171875 -0.421875 C -3.792969 -0.421875 -4.355469 -0.527344 -4.851563 -0.746094 C -5.34375 -0.960938 -5.71875 -1.277344 -5.976563 -1.691406 C -6.234375 -2.101563 -6.363281 -2.554688 -6.363281 -3.046875 C -6.363281 -3.816406 -6.039063 -4.421875 -5.390625 -4.863281 L -6.222656 -4.863281 L -6.222656 -5.8125 L 2.386719 -5.8125 Z M -3.128906 -1.507813 C -2.328125 -1.503906 -1.726563 -1.671875 -1.328125 -2.011719 C -0.925781 -2.34375 -0.726563 -2.746094 -0.726563 -3.21875 C -0.726563 -3.664063 -0.914063 -4.050781 -1.296875 -4.375 C -1.671875 -4.699219 -2.253906 -4.863281 -3.035156 -4.863281 C -3.863281 -4.863281 -4.484375 -4.691406 -4.902344 -4.351563 C -5.320313 -4.007813 -5.53125 -3.605469 -5.53125 -3.148438 C -5.53125 -2.6875 -5.335938 -2.300781 -4.949219 -1.984375 C -4.558594 -1.664063 -3.953125 -1.503906 -3.128906 -1.507813 Z M -3.128906 -1.507813 "/>
</symbol>
<symbol overflow="visible" id="glyph2-5">
<path style="stroke:none;" d="M 0 -4.867188 L -0.914063 -4.867188 C -0.210938 -4.378906 0.140625 -3.722656 0.140625 -2.894531 C 0.140625 -2.527344 0.0703125 -2.183594 -0.0703125 -1.867188 C -0.210938 -1.546875 -0.386719 -1.308594 -0.597656 -1.15625 C -0.808594 -1 -1.070313 -0.894531 -1.382813 -0.832031 C -1.589844 -0.789063 -1.917969 -0.765625 -2.367188 -0.769531 L -6.222656 -0.769531 L -6.222656 -1.824219 L -2.773438 -1.824219 C -2.21875 -1.820313 -1.847656 -1.84375 -1.65625 -1.886719 C -1.378906 -1.949219 -1.160156 -2.089844 -1.003906 -2.308594 C -0.839844 -2.523438 -0.761719 -2.789063 -0.765625 -3.105469 C -0.761719 -3.417969 -0.84375 -3.714844 -1.007813 -3.996094 C -1.171875 -4.273438 -1.390625 -4.46875 -1.671875 -4.585938 C -1.945313 -4.699219 -2.351563 -4.757813 -2.886719 -4.757813 L -6.222656 -4.757813 L -6.222656 -5.8125 L 0 -5.8125 Z M 0 -4.867188 "/>
</symbol>
<symbol overflow="visible" id="glyph2-6">
<path style="stroke:none;" d="M 0 -0.789063 L -6.222656 -0.792969 L -6.222656 -1.742188 L -5.335938 -1.742188 C -6.019531 -2.195313 -6.363281 -2.855469 -6.363281 -3.722656 C -6.363281 -4.089844 -6.292969 -4.433594 -6.160156 -4.753906 C -6.023438 -5.066406 -5.847656 -5.304688 -5.632813 -5.460938 C -5.410156 -5.617188 -5.152344 -5.726563 -4.851563 -5.789063 C -4.65625 -5.828125 -4.3125 -5.847656 -3.824219 -5.847656 L 0 -5.847656 L 0 -4.792969 L -3.785156 -4.792969 C -4.214844 -4.792969 -4.535156 -4.75 -4.75 -4.667969 C -4.960938 -4.585938 -5.128906 -4.441406 -5.257813 -4.234375 C -5.382813 -4.023438 -5.449219 -3.777344 -5.449219 -3.5 C -5.449219 -3.046875 -5.304688 -2.660156 -5.019531 -2.335938 C -4.734375 -2.007813 -4.195313 -1.84375 -3.398438 -1.847656 L 0 -1.84375 Z M 0 -0.789063 "/>
</symbol>
<symbol overflow="visible" id="glyph2-7">
<path style="stroke:none;" d="M -2.277344 -4.851563 L -2.144531 -5.890625 C -1.425781 -5.773438 -0.863281 -5.484375 -0.464844 -5.019531 C -0.0585938 -4.550781 0.140625 -3.976563 0.140625 -3.296875 C 0.140625 -2.445313 -0.136719 -1.761719 -0.695313 -1.246094 C -1.25 -0.726563 -2.046875 -0.46875 -3.085938 -0.46875 C -3.753906 -0.46875 -4.34375 -0.578125 -4.851563 -0.800781 C -5.355469 -1.023438 -5.730469 -1.363281 -5.984375 -1.820313 C -6.234375 -2.273438 -6.363281 -2.769531 -6.363281 -3.304688 C -6.363281 -3.980469 -6.191406 -4.53125 -5.847656 -4.964844 C -5.503906 -5.390625 -5.019531 -5.667969 -4.394531 -5.789063 L -4.234375 -4.765625 C -4.652344 -4.664063 -4.96875 -4.492188 -5.179688 -4.246094 C -5.390625 -3.996094 -5.496094 -3.695313 -5.496094 -3.347656 C -5.496094 -2.8125 -5.304688 -2.382813 -4.921875 -2.050781 C -4.539063 -1.71875 -3.9375 -1.550781 -3.117188 -1.554688 C -2.28125 -1.550781 -1.671875 -1.710938 -1.292969 -2.035156 C -0.914063 -2.351563 -0.726563 -2.769531 -0.726563 -3.289063 C -0.726563 -3.695313 -0.851563 -4.042969 -1.105469 -4.324219 C -1.359375 -4.601563 -1.75 -4.777344 -2.277344 -4.851563 Z M -2.277344 -4.851563 "/>
</symbol>
<symbol overflow="visible" id="glyph2-8">
<path style="stroke:none;" d="M 2.398438 -0.742188 L 1.40625 -0.625 C 1.46875 -0.855469 1.5 -1.058594 1.5 -1.230469 C 1.5 -1.464844 1.460938 -1.652344 1.382813 -1.792969 C 1.304688 -1.933594 1.195313 -2.046875 1.054688 -2.140625 C 0.949219 -2.203125 0.6875 -2.3125 0.269531 -2.460938 C 0.210938 -2.480469 0.125 -2.511719 0.0117188 -2.554688 L -6.222656 -0.195313 L -6.222656 -1.332031 L -2.617188 -2.625 C -2.160156 -2.789063 -1.679688 -2.9375 -1.175781 -3.078125 C -1.65625 -3.195313 -2.128906 -3.339844 -2.59375 -3.507813 L -6.222656 -4.839844 L -6.222656 -5.894531 L 0.105469 -3.527344 C 0.789063 -3.273438 1.257813 -3.074219 1.519531 -2.9375 C 1.863281 -2.746094 2.117188 -2.53125 2.28125 -2.289063 C 2.4375 -2.042969 2.519531 -1.753906 2.523438 -1.421875 C 2.519531 -1.214844 2.476563 -0.988281 2.398438 -0.742188 Z M 2.398438 -0.742188 "/>
</symbol>
<symbol overflow="visible" id="glyph2-9">
<path style="stroke:none;" d="M -4.234375 -0.5 C -5.246094 -0.496094 -6.0625 -0.601563 -6.6875 -0.8125 C -7.304688 -1.019531 -7.785156 -1.328125 -8.121094 -1.742188 C -8.457031 -2.152344 -8.625 -2.671875 -8.625 -3.300781 C -8.625 -3.757813 -8.53125 -4.164063 -8.347656 -4.511719 C -8.160156 -4.859375 -7.890625 -5.144531 -7.542969 -5.371094 C -7.191406 -5.59375 -6.765625 -5.773438 -6.265625 -5.90625 C -5.761719 -6.035156 -5.085938 -6.097656 -4.234375 -6.101563 C -3.222656 -6.097656 -2.410156 -5.996094 -1.792969 -5.789063 C -1.175781 -5.578125 -0.695313 -5.265625 -0.359375 -4.859375 C -0.0195313 -4.445313 0.144531 -3.925781 0.148438 -3.296875 C 0.144531 -2.464844 -0.148438 -1.816406 -0.742188 -1.347656 C -1.457031 -0.78125 -2.621094 -0.496094 -4.234375 -0.5 Z M -4.234375 -1.582031 C -2.824219 -1.582031 -1.886719 -1.746094 -1.417969 -2.074219 C -0.949219 -2.402344 -0.714844 -2.808594 -0.71875 -3.296875 C -0.714844 -3.777344 -0.949219 -4.183594 -1.421875 -4.519531 C -1.886719 -4.847656 -2.824219 -5.015625 -4.234375 -5.015625 C -5.648438 -5.015625 -6.589844 -4.847656 -7.054688 -4.519531 C -7.515625 -4.1875 -7.746094 -3.777344 -7.75 -3.289063 C -7.746094 -2.800781 -7.542969 -2.414063 -7.136719 -2.128906 C -6.613281 -1.761719 -5.644531 -1.582031 -4.234375 -1.582031 Z M -4.234375 -1.582031 "/>
</symbol>
<symbol overflow="visible" id="glyph2-10">
<path style="stroke:none;" d="M 0 -1.089844 L -1.203125 -1.089844 L -1.199219 -2.289063 L 0 -2.289063 Z M 0 -1.089844 "/>
</symbol>
<symbol overflow="visible" id="glyph2-11">
<path style="stroke:none;" d="M -1.011719 -6.039063 L 0 -6.039063 L 0 -0.363281 C -0.253906 -0.355469 -0.496094 -0.394531 -0.734375 -0.488281 C -1.117188 -0.628906 -1.5 -0.859375 -1.875 -1.179688 C -2.25 -1.496094 -2.683594 -1.957031 -3.175781 -2.5625 C -3.941406 -3.492188 -4.546875 -4.125 -4.992188 -4.453125 C -5.4375 -4.78125 -5.859375 -4.945313 -6.265625 -4.945313 C -6.679688 -4.945313 -7.03125 -4.792969 -7.320313 -4.496094 C -7.601563 -4.195313 -7.746094 -3.808594 -7.75 -3.328125 C -7.746094 -2.820313 -7.59375 -2.414063 -7.292969 -2.109375 C -6.984375 -1.804688 -6.5625 -1.648438 -6.03125 -1.648438 L -6.140625 -0.5625 C -6.945313 -0.636719 -7.558594 -0.914063 -7.988281 -1.402344 C -8.410156 -1.882813 -8.625 -2.535156 -8.625 -3.351563 C -8.625 -4.175781 -8.394531 -4.828125 -7.9375 -5.308594 C -7.480469 -5.789063 -6.914063 -6.027344 -6.242188 -6.03125 C -5.894531 -6.027344 -5.558594 -5.957031 -5.226563 -5.820313 C -4.890625 -5.675781 -4.539063 -5.441406 -4.175781 -5.117188 C -3.804688 -4.789063 -3.300781 -4.25 -2.664063 -3.492188 C -2.128906 -2.859375 -1.769531 -2.453125 -1.582031 -2.273438 C -1.394531 -2.09375 -1.203125 -1.945313 -1.011719 -1.828125 Z M -1.011719 -6.039063 "/>
</symbol>
<symbol overflow="visible" id="glyph2-12">
<path style="stroke:none;" d="M 0 -3.878906 L -2.054688 -3.878906 L -2.054688 -0.152344 L -3.023438 -0.152344 L -8.589844 -4.074219 L -8.589844 -4.933594 L -3.023438 -4.933594 L -3.023438 -6.09375 L -2.054688 -6.09375 L -2.054688 -4.933594 L 0 -4.933594 Z M -3.023438 -3.878906 L -6.898438 -3.878906 L -3.023438 -1.191406 Z M -3.023438 -3.878906 "/>
</symbol>
<symbol overflow="visible" id="glyph2-13">
<path style="stroke:none;" d="M -6.484375 -5.96875 L -6.40625 -4.921875 C -6.8125 -4.828125 -7.113281 -4.695313 -7.304688 -4.523438 C -7.605469 -4.238281 -7.757813 -3.886719 -7.757813 -3.46875 C -7.757813 -3.132813 -7.664063 -2.835938 -7.476563 -2.585938 C -7.234375 -2.25 -6.878906 -1.988281 -6.414063 -1.796875 C -5.949219 -1.605469 -5.289063 -1.507813 -4.429688 -1.5 C -4.8125 -1.753906 -5.097656 -2.0625 -5.289063 -2.433594 C -5.472656 -2.796875 -5.566406 -3.183594 -5.570313 -3.585938 C -5.566406 -4.289063 -5.308594 -4.886719 -4.792969 -5.382813 C -4.277344 -5.875 -3.609375 -6.121094 -2.789063 -6.125 C -2.25 -6.121094 -1.746094 -6.003906 -1.285156 -5.773438 C -0.816406 -5.539063 -0.460938 -5.222656 -0.21875 -4.816406 C 0.0273438 -4.410156 0.144531 -3.949219 0.148438 -3.433594 C 0.144531 -2.554688 -0.175781 -1.835938 -0.820313 -1.285156 C -1.46875 -0.726563 -2.535156 -0.449219 -4.019531 -0.453125 C -5.675781 -0.449219 -6.882813 -0.757813 -7.640625 -1.371094 C -8.296875 -1.90625 -8.625 -2.625 -8.625 -3.535156 C -8.625 -4.207031 -8.433594 -4.761719 -8.054688 -5.195313 C -7.675781 -5.625 -7.152344 -5.882813 -6.484375 -5.96875 Z M -2.78125 -1.664063 C -2.417969 -1.664063 -2.070313 -1.738281 -1.738281 -1.894531 C -1.40625 -2.042969 -1.152344 -2.261719 -0.980469 -2.542969 C -0.800781 -2.820313 -0.714844 -3.109375 -0.71875 -3.414063 C -0.714844 -3.859375 -0.894531 -4.242188 -1.257813 -4.566406 C -1.613281 -4.882813 -2.101563 -5.042969 -2.722656 -5.046875 C -3.3125 -5.042969 -3.78125 -4.886719 -4.125 -4.570313 C -4.46875 -4.25 -4.640625 -3.851563 -4.640625 -3.375 C -4.640625 -2.898438 -4.46875 -2.492188 -4.128906 -2.160156 C -3.785156 -1.828125 -3.335938 -1.664063 -2.78125 -1.664063 Z M -2.78125 -1.664063 "/>
</symbol>
<symbol overflow="visible" id="glyph2-14">
<path style="stroke:none;" d="M -4.65625 -2.121094 C -4.816406 -1.683594 -5.046875 -1.359375 -5.34375 -1.148438 C -5.640625 -0.9375 -5.996094 -0.832031 -6.410156 -0.832031 C -7.035156 -0.832031 -7.558594 -1.054688 -7.984375 -1.503906 C -8.410156 -1.953125 -8.625 -2.550781 -8.625 -3.300781 C -8.625 -4.046875 -8.40625 -4.652344 -7.972656 -5.109375 C -7.535156 -5.566406 -7.003906 -5.792969 -6.382813 -5.796875 C -5.976563 -5.792969 -5.628906 -5.6875 -5.339844 -5.480469 C -5.042969 -5.269531 -4.816406 -4.953125 -4.65625 -4.53125 C -4.480469 -5.054688 -4.203125 -5.457031 -3.824219 -5.734375 C -3.4375 -6.007813 -2.980469 -6.144531 -2.453125 -6.148438 C -1.714844 -6.144531 -1.097656 -5.886719 -0.601563 -5.367188 C -0.101563 -4.84375 0.144531 -4.160156 0.148438 -3.316406 C 0.144531 -2.46875 -0.101563 -1.785156 -0.605469 -1.265625 C -1.105469 -0.746094 -1.734375 -0.484375 -2.484375 -0.488281 C -3.039063 -0.484375 -3.503906 -0.625 -3.886719 -0.910156 C -4.261719 -1.191406 -4.519531 -1.597656 -4.65625 -2.121094 Z M -6.445313 -1.910156 C -6.039063 -1.910156 -5.707031 -2.039063 -5.449219 -2.300781 C -5.191406 -2.5625 -5.0625 -2.902344 -5.0625 -3.324219 C -5.0625 -3.726563 -5.1875 -4.058594 -5.445313 -4.320313 C -5.695313 -4.578125 -6.011719 -4.710938 -6.386719 -4.710938 C -6.773438 -4.710938 -7.097656 -4.574219 -7.363281 -4.308594 C -7.625 -4.039063 -7.757813 -3.707031 -7.757813 -3.3125 C -7.757813 -2.90625 -7.628906 -2.574219 -7.371094 -2.308594 C -7.113281 -2.042969 -6.804688 -1.910156 -6.445313 -1.910156 Z M -2.476563 -1.570313 C -2.175781 -1.570313 -1.886719 -1.640625 -1.605469 -1.785156 C -1.324219 -1.925781 -1.105469 -2.136719 -0.949219 -2.421875 C -0.792969 -2.699219 -0.714844 -3.003906 -0.71875 -3.328125 C -0.714844 -3.832031 -0.875 -4.246094 -1.203125 -4.578125 C -1.523438 -4.902344 -1.9375 -5.066406 -2.441406 -5.070313 C -2.945313 -5.066406 -3.367188 -4.898438 -3.703125 -4.5625 C -4.035156 -4.222656 -4.199219 -3.800781 -4.203125 -3.292969 C -4.199219 -2.796875 -4.035156 -2.382813 -3.710938 -2.058594 C -3.378906 -1.730469 -2.96875 -1.570313 -2.476563 -1.570313 Z M -2.476563 -1.570313 "/>
</symbol>
<symbol overflow="visible" id="glyph2-15">
<path style="stroke:none;" d="M 0 -4.46875 L 0 -3.414063 L -6.71875 -3.417969 C -6.476563 -3.160156 -6.234375 -2.828125 -5.996094 -2.417969 C -5.75 -2.003906 -5.570313 -1.632813 -5.449219 -1.308594 L -6.46875 -1.308594 C -6.742188 -1.894531 -7.078125 -2.410156 -7.476563 -2.851563 C -7.871094 -3.292969 -8.253906 -3.605469 -8.625 -3.792969 L -8.625 -4.472656 Z M 0 -4.46875 "/>
</symbol>
</g>
</defs>
<g id="surface31">
<rect x="0" y="0" width="504" height="504" style="fill:rgb(100%,100%,100%);fill-opacity:1;stroke:none;"/>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph0-1" x="250.398438" y="34.675781"/>
  <use xlink:href="#glyph0-2" x="260.797656" y="34.675781"/>
  <use xlink:href="#glyph0-3" x="269.59375" y="34.675781"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph1-1" x="135.996094" y="485.28125"/>
  <use xlink:href="#glyph1-2" x="144" y="485.28125"/>
  <use xlink:href="#glyph1-3" x="150" y="485.28125"/>
  <use xlink:href="#glyph1-4" x="156.673828" y="485.28125"/>
  <use xlink:href="#glyph1-5" x="160.669922" y="485.28125"/>
  <use xlink:href="#glyph1-6" x="167.34375" y="485.28125"/>
  <use xlink:href="#glyph1-3" x="174.017578" y="485.28125"/>
  <use xlink:href="#glyph1-7" x="180.691406" y="485.28125"/>
  <use xlink:href="#glyph1-8" x="187.365234" y="485.28125"/>
  <use xlink:href="#glyph1-9" x="196.03125" y="485.28125"/>
  <use xlink:href="#glyph1-10" x="202.705078" y="485.28125"/>
  <use xlink:href="#glyph1-11" x="212.701172" y="485.28125"/>
  <use xlink:href="#glyph1-3" x="219.375" y="485.28125"/>
  <use xlink:href="#glyph1-4" x="226.048828" y="485.28125"/>
  <use xlink:href="#glyph1-7" x="230.044922" y="485.28125"/>
  <use xlink:href="#glyph1-12" x="236.71875" y="485.28125"/>
  <use xlink:href="#glyph1-13" x="246.052734" y="485.28125"/>
  <use xlink:href="#glyph1-7" x="249.386719" y="485.28125"/>
  <use xlink:href="#glyph1-14" x="256.060547" y="485.28125"/>
  <use xlink:href="#glyph1-15" x="264.726563" y="485.28125"/>
  <use xlink:href="#glyph1-16" x="271.400391" y="485.28125"/>
  <use xlink:href="#glyph1-17" x="274.066406" y="485.28125"/>
  <use xlink:href="#glyph1-18" x="276.732422" y="485.28125"/>
  <use xlink:href="#glyph1-4" x="283.40625" y="485.28125"/>
  <use xlink:href="#glyph1-3" x="287.402344" y="485.28125"/>
  <use xlink:href="#glyph1-19" x="294.076172" y="485.28125"/>
  <use xlink:href="#glyph1-7" x="300.75" y="485.28125"/>
  <use xlink:href="#glyph1-20" x="307.423828" y="485.28125"/>
  <use xlink:href="#glyph1-3" x="315.427734" y="485.28125"/>
  <use xlink:href="#glyph1-4" x="322.101563" y="485.28125"/>
  <use xlink:href="#glyph1-7" x="326.097656" y="485.28125"/>
  <use xlink:href="#glyph1-21" x="332.771484" y="485.28125"/>
  <use xlink:href="#glyph1-5" x="340.775391" y="485.28125"/>
  <use xlink:href="#glyph1-22" x="347.449219" y="485.28125"/>
  <use xlink:href="#glyph1-3" x="353.449219" y="485.28125"/>
  <use xlink:href="#glyph1-7" x="360.123047" y="485.28125"/>
  <use xlink:href="#glyph1-14" x="366.796875" y="485.28125"/>
  <use xlink:href="#glyph1-17" x="375.462891" y="485.28125"/>
  <use xlink:href="#glyph1-5" x="378.128906" y="485.28125"/>
  <use xlink:href="#glyph1-22" x="384.802734" y="485.28125"/>
  <use xlink:href="#glyph1-22" x="390.802734" y="485.28125"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-1" x="12.960938" y="273.148438"/>
  <use xlink:href="#glyph2-2" x="12.960938" y="265.818359"/>
  <use xlink:href="#glyph2-3" x="12.960938" y="261.822266"/>
  <use xlink:href="#glyph2-4" x="12.960938" y="255.148438"/>
  <use xlink:href="#glyph2-5" x="12.960938" y="248.474609"/>
  <use xlink:href="#glyph2-3" x="12.960938" y="241.800781"/>
  <use xlink:href="#glyph2-6" x="12.960938" y="235.126953"/>
  <use xlink:href="#glyph2-7" x="12.960938" y="228.453125"/>
  <use xlink:href="#glyph2-8" x="12.960938" y="222.453125"/>
</g>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 74.398438 430.558594 L 458.398438 430.558594 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 74.398438 430.558594 L 74.398438 437.761719 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 151.199219 430.558594 L 151.199219 437.761719 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 228 430.558594 L 228 437.761719 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 304.800781 430.558594 L 304.800781 437.761719 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 381.601563 430.558594 L 381.601563 437.761719 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 458.398438 430.558594 L 458.398438 437.761719 "/>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph1-23" x="66.058594" y="456.480469"/>
  <use xlink:href="#glyph1-24" x="72.732422" y="456.480469"/>
  <use xlink:href="#glyph1-25" x="76.066406" y="456.480469"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph1-23" x="142.859375" y="456.480469"/>
  <use xlink:href="#glyph1-24" x="149.533203" y="456.480469"/>
  <use xlink:href="#glyph1-26" x="152.867188" y="456.480469"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph1-23" x="219.660156" y="456.480469"/>
  <use xlink:href="#glyph1-24" x="226.333984" y="456.480469"/>
  <use xlink:href="#glyph1-27" x="229.667969" y="456.480469"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph1-23" x="296.460938" y="456.480469"/>
  <use xlink:href="#glyph1-24" x="303.134766" y="456.480469"/>
  <use xlink:href="#glyph1-28" x="306.46875" y="456.480469"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph1-23" x="373.261719" y="456.480469"/>
  <use xlink:href="#glyph1-24" x="379.935547" y="456.480469"/>
  <use xlink:href="#glyph1-29" x="383.269531" y="456.480469"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph1-30" x="450.058594" y="456.480469"/>
  <use xlink:href="#glyph1-24" x="456.732422" y="456.480469"/>
  <use xlink:href="#glyph1-23" x="460.066406" y="456.480469"/>
</g>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 59.039063 416.800781 L 59.039063 72.800781 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 59.039063 416.800781 L 51.839844 416.800781 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 59.039063 348 L 51.839844 348 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 59.039063 279.199219 L 51.839844 279.199219 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 59.039063 210.398438 L 51.839844 210.398438 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 59.039063 141.601563 L 51.839844 141.601563 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 59.039063 72.800781 L 51.839844 72.800781 "/>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-9" x="41.761719" y="425.140625"/>
  <use xlink:href="#glyph2-10" x="41.761719" y="418.466797"/>
  <use xlink:href="#glyph2-9" x="41.761719" y="415.132813"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-9" x="41.761719" y="356.339844"/>
  <use xlink:href="#glyph2-10" x="41.761719" y="349.666016"/>
  <use xlink:href="#glyph2-11" x="41.761719" y="346.332031"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-9" x="41.761719" y="287.539063"/>
  <use xlink:href="#glyph2-10" x="41.761719" y="280.865234"/>
  <use xlink:href="#glyph2-12" x="41.761719" y="277.53125"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-9" x="41.761719" y="218.738281"/>
  <use xlink:href="#glyph2-10" x="41.761719" y="212.064453"/>
  <use xlink:href="#glyph2-13" x="41.761719" y="208.730469"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-9" x="41.761719" y="149.941406"/>
  <use xlink:href="#glyph2-10" x="41.761719" y="143.267578"/>
  <use xlink:href="#glyph2-14" x="41.761719" y="139.933594"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-15" x="41.761719" y="81.140625"/>
  <use xlink:href="#glyph2-10" x="41.761719" y="74.466797"/>
  <use xlink:href="#glyph2-9" x="41.761719" y="71.132813"/>
</g>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 74.398438 416.800781 L 458.398438 416.800781 L 458.398438 72.800781 L 74.398438 72.800781 Z M 74.398438 416.800781 "/>
</g>
</svg>
