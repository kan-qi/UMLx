<?xml version="1.0" encoding="UTF-8"?>
<svg xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" width="360pt" height="360pt" viewBox="0 0 360 360" version="1.1">
<defs>
<g>
<symbol overflow="visible" id="glyph0-0">
<path style="stroke:none;" d="M 1.5 0 L 1.5 -7.5 L 7.5 -7.5 L 7.5 0 Z M 1.6875 -0.1875 L 7.3125 -0.1875 L 7.3125 -7.3125 L 1.6875 -7.3125 Z M 1.6875 -0.1875 "/>
</symbol>
<symbol overflow="visible" id="glyph0-1">
<path style="stroke:none;" d="M 6.039063 -1.015625 L 6.039063 0 L 0.363281 0 C 0.355469 -0.253906 0.394531 -0.496094 0.484375 -0.734375 C 0.628906 -1.117188 0.859375 -1.5 1.179688 -1.875 C 1.492188 -2.25 1.953125 -2.683594 2.5625 -3.175781 C 3.492188 -3.941406 4.125 -4.546875 4.453125 -4.992188 C 4.78125 -5.4375 4.945313 -5.859375 4.945313 -6.265625 C 4.945313 -6.679688 4.792969 -7.03125 4.496094 -7.320313 C 4.191406 -7.601563 3.804688 -7.746094 3.328125 -7.75 C 2.820313 -7.746094 2.414063 -7.59375 2.109375 -7.292969 C 1.804688 -6.984375 1.648438 -6.5625 1.648438 -6.03125 L 0.5625 -6.140625 C 0.632813 -6.945313 0.910156 -7.558594 1.398438 -7.988281 C 1.878906 -8.410156 2.53125 -8.625 3.351563 -8.625 C 4.171875 -8.625 4.824219 -8.394531 5.308594 -7.9375 C 5.789063 -7.480469 6.027344 -6.914063 6.03125 -6.242188 C 6.027344 -5.894531 5.957031 -5.558594 5.820313 -5.226563 C 5.675781 -4.890625 5.441406 -4.539063 5.117188 -4.175781 C 4.789063 -3.804688 4.25 -3.300781 3.492188 -2.664063 C 2.859375 -2.128906 2.453125 -1.769531 2.273438 -1.582031 C 2.09375 -1.394531 1.945313 -1.203125 1.828125 -1.015625 Z M 6.039063 -1.015625 "/>
</symbol>
<symbol overflow="visible" id="glyph0-2">
<path style="stroke:none;" d="M 0.5 -2.25 L 1.605469 -2.34375 C 1.683594 -1.804688 1.871094 -1.398438 2.175781 -1.125 C 2.472656 -0.851563 2.835938 -0.714844 3.257813 -0.71875 C 3.765625 -0.714844 4.195313 -0.90625 4.546875 -1.292969 C 4.898438 -1.671875 5.074219 -2.179688 5.074219 -2.820313 C 5.074219 -3.414063 4.902344 -3.890625 4.566406 -4.242188 C 4.226563 -4.589844 3.785156 -4.761719 3.242188 -4.765625 C 2.898438 -4.761719 2.59375 -4.683594 2.320313 -4.53125 C 2.046875 -4.375 1.832031 -4.175781 1.675781 -3.929688 L 0.6875 -4.0625 L 1.515625 -8.472656 L 5.789063 -8.472656 L 5.789063 -7.464844 L 2.359375 -7.464844 L 1.898438 -5.15625 C 2.414063 -5.515625 2.953125 -5.695313 3.523438 -5.695313 C 4.269531 -5.695313 4.902344 -5.433594 5.421875 -4.914063 C 5.933594 -4.394531 6.191406 -3.726563 6.195313 -2.914063 C 6.191406 -2.132813 5.964844 -1.460938 5.515625 -0.898438 C 4.960938 -0.199219 4.210938 0.144531 3.257813 0.148438 C 2.476563 0.144531 1.835938 -0.0703125 1.34375 -0.507813 C 0.84375 -0.941406 0.5625 -1.523438 0.5 -2.25 Z M 0.5 -2.25 "/>
</symbol>
<symbol overflow="visible" id="glyph0-3">
<path style="stroke:none;" d="M 0.695313 -6.527344 C 0.691406 -7.136719 0.847656 -7.65625 1.160156 -8.089844 C 1.46875 -8.515625 1.914063 -8.730469 2.5 -8.734375 C 3.039063 -8.730469 3.484375 -8.539063 3.839844 -8.15625 C 4.191406 -7.773438 4.371094 -7.207031 4.371094 -6.460938 C 4.371094 -5.734375 4.191406 -5.175781 3.832031 -4.785156 C 3.472656 -4.390625 3.03125 -4.195313 2.515625 -4.195313 C 1.992188 -4.195313 1.558594 -4.386719 1.214844 -4.773438 C 0.863281 -5.160156 0.691406 -5.746094 0.695313 -6.527344 Z M 2.53125 -8.007813 C 2.269531 -8.003906 2.050781 -7.890625 1.878906 -7.667969 C 1.703125 -7.4375 1.617188 -7.023438 1.617188 -6.421875 C 1.617188 -5.867188 1.703125 -5.476563 1.878906 -5.257813 C 2.054688 -5.03125 2.273438 -4.921875 2.53125 -4.921875 C 2.796875 -4.921875 3.015625 -5.035156 3.191406 -5.261719 C 3.363281 -5.488281 3.449219 -5.902344 3.453125 -6.503906 C 3.449219 -7.058594 3.363281 -7.445313 3.1875 -7.671875 C 3.007813 -7.890625 2.789063 -8.003906 2.53125 -8.007813 Z M 2.539063 0.316406 L 7.234375 -8.734375 L 8.09375 -8.734375 L 3.410156 0.316406 Z M 6.25 -2.015625 C 6.246094 -2.632813 6.402344 -3.152344 6.714844 -3.582031 C 7.023438 -4.007813 7.472656 -4.222656 8.0625 -4.226563 C 8.601563 -4.222656 9.046875 -4.03125 9.398438 -3.648438 C 9.75 -3.261719 9.925781 -2.695313 9.929688 -1.953125 C 9.925781 -1.21875 9.746094 -0.660156 9.394531 -0.269531 C 9.035156 0.121094 8.59375 0.316406 8.070313 0.316406 C 7.546875 0.316406 7.113281 0.125 6.769531 -0.265625 C 6.417969 -0.652344 6.246094 -1.238281 6.25 -2.015625 Z M 8.09375 -3.5 C 7.824219 -3.496094 7.605469 -3.382813 7.433594 -3.160156 C 7.257813 -2.929688 7.171875 -2.515625 7.171875 -1.910156 C 7.171875 -1.363281 7.257813 -0.976563 7.433594 -0.75 C 7.609375 -0.523438 7.828125 -0.410156 8.085938 -0.410156 C 8.355469 -0.410156 8.574219 -0.523438 8.75 -0.75 C 8.921875 -0.976563 9.011719 -1.390625 9.011719 -1.992188 C 9.011719 -2.546875 8.921875 -2.933594 8.746094 -3.160156 C 8.570313 -3.382813 8.351563 -3.496094 8.09375 -3.5 Z M 8.09375 -3.5 "/>
</symbol>
<symbol overflow="visible" id="glyph0-4">
<path style="stroke:none;" d="M 0.5 -4.234375 C 0.496094 -5.246094 0.601563 -6.0625 0.8125 -6.6875 C 1.019531 -7.304688 1.328125 -7.785156 1.742188 -8.121094 C 2.148438 -8.457031 2.667969 -8.625 3.296875 -8.625 C 3.757813 -8.625 4.164063 -8.53125 4.511719 -8.347656 C 4.855469 -8.160156 5.140625 -7.890625 5.371094 -7.542969 C 5.59375 -7.191406 5.773438 -6.765625 5.90625 -6.265625 C 6.035156 -5.761719 6.097656 -5.085938 6.101563 -4.234375 C 6.097656 -3.226563 5.996094 -2.414063 5.789063 -1.796875 C 5.578125 -1.175781 5.265625 -0.695313 4.859375 -0.359375 C 4.445313 -0.0195313 3.925781 0.144531 3.296875 0.148438 C 2.464844 0.144531 1.816406 -0.148438 1.347656 -0.742188 C 0.78125 -1.457031 0.496094 -2.621094 0.5 -4.234375 Z M 1.582031 -4.234375 C 1.582031 -2.824219 1.746094 -1.886719 2.074219 -1.417969 C 2.402344 -0.949219 2.808594 -0.714844 3.296875 -0.71875 C 3.777344 -0.714844 4.183594 -0.949219 4.519531 -1.421875 C 4.847656 -1.886719 5.015625 -2.824219 5.015625 -4.234375 C 5.015625 -5.648438 4.847656 -6.589844 4.519531 -7.054688 C 4.183594 -7.515625 3.773438 -7.746094 3.289063 -7.75 C 2.800781 -7.746094 2.414063 -7.542969 2.125 -7.136719 C 1.761719 -6.613281 1.582031 -5.644531 1.582031 -4.234375 Z M 1.582031 -4.234375 "/>
</symbol>
<symbol overflow="visible" id="glyph1-0">
<path style="stroke:none;" d="M 1.800781 0 L 1.800781 -9 L 9 -9 L 9 0 Z M 2.023438 -0.226563 L 8.773438 -0.226563 L 8.773438 -8.773438 L 2.023438 -8.773438 Z M 2.023438 -0.226563 "/>
</symbol>
<symbol overflow="visible" id="glyph1-1">
<path style="stroke:none;" d="M 1.039063 -10.308594 L 4.84375 -10.308594 C 5.699219 -10.304688 6.351563 -10.238281 6.804688 -10.109375 C 7.40625 -9.929688 7.925781 -9.613281 8.359375 -9.160156 C 8.789063 -8.703125 9.117188 -8.148438 9.34375 -7.492188 C 9.566406 -6.832031 9.679688 -6.019531 9.683594 -5.054688 C 9.679688 -4.203125 9.574219 -3.472656 9.367188 -2.863281 C 9.105469 -2.109375 8.738281 -1.5 8.261719 -1.039063 C 7.898438 -0.683594 7.410156 -0.410156 6.800781 -0.21875 C 6.335938 -0.0703125 5.722656 0 4.957031 0 L 1.039063 0 Z M 3.121094 -8.5625 L 3.121094 -1.738281 L 4.675781 -1.738281 C 5.253906 -1.734375 5.671875 -1.765625 5.933594 -1.835938 C 6.269531 -1.914063 6.550781 -2.058594 6.773438 -2.261719 C 6.996094 -2.464844 7.175781 -2.796875 7.320313 -3.257813 C 7.457031 -3.71875 7.527344 -4.347656 7.53125 -5.148438 C 7.527344 -5.941406 7.457031 -6.550781 7.320313 -6.980469 C 7.175781 -7.402344 6.980469 -7.738281 6.726563 -7.980469 C 6.472656 -8.21875 6.152344 -8.378906 5.765625 -8.464844 C 5.472656 -8.527344 4.902344 -8.558594 4.058594 -8.5625 Z M 3.121094 -8.5625 "/>
</symbol>
<symbol overflow="visible" id="glyph1-2">
<path style="stroke:none;" d="M 1.035156 -8.480469 L 1.035156 -10.308594 L 3.007813 -10.308594 L 3.007813 -8.480469 Z M 1.035156 0 L 1.035156 -7.46875 L 3.007813 -7.46875 L 3.007813 0 Z M 1.035156 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-3">
<path style="stroke:none;" d="M 0.335938 -2.128906 L 2.320313 -2.433594 C 2.402344 -2.042969 2.570313 -1.75 2.832031 -1.554688 C 3.085938 -1.351563 3.449219 -1.253906 3.917969 -1.257813 C 4.425781 -1.253906 4.808594 -1.347656 5.070313 -1.539063 C 5.238281 -1.667969 5.324219 -1.84375 5.328125 -2.066406 C 5.324219 -2.214844 5.277344 -2.339844 5.1875 -2.441406 C 5.085938 -2.53125 4.867188 -2.617188 4.527344 -2.699219 C 2.929688 -3.046875 1.917969 -3.367188 1.496094 -3.664063 C 0.902344 -4.0625 0.609375 -4.625 0.613281 -5.34375 C 0.609375 -5.988281 0.863281 -6.53125 1.378906 -6.972656 C 1.886719 -7.414063 2.679688 -7.632813 3.753906 -7.636719 C 4.773438 -7.632813 5.53125 -7.46875 6.03125 -7.136719 C 6.523438 -6.800781 6.867188 -6.308594 7.058594 -5.660156 L 5.195313 -5.316406 C 5.113281 -5.601563 4.960938 -5.824219 4.742188 -5.980469 C 4.515625 -6.132813 4.199219 -6.210938 3.789063 -6.214844 C 3.265625 -6.210938 2.894531 -6.136719 2.671875 -5.996094 C 2.519531 -5.890625 2.441406 -5.757813 2.445313 -5.597656 C 2.441406 -5.453125 2.507813 -5.335938 2.644531 -5.238281 C 2.816406 -5.105469 3.433594 -4.917969 4.488281 -4.683594 C 5.539063 -4.441406 6.273438 -4.148438 6.695313 -3.804688 C 7.105469 -3.449219 7.3125 -2.960938 7.3125 -2.335938 C 7.3125 -1.648438 7.023438 -1.058594 6.453125 -0.570313 C 5.878906 -0.078125 5.035156 0.164063 3.917969 0.167969 C 2.898438 0.164063 2.09375 -0.0390625 1.5 -0.449219 C 0.90625 -0.859375 0.515625 -1.417969 0.335938 -2.128906 Z M 0.335938 -2.128906 "/>
</symbol>
<symbol overflow="visible" id="glyph1-4">
<path style="stroke:none;" d="M 4.457031 -7.46875 L 4.457031 -5.890625 L 3.109375 -5.890625 L 3.109375 -2.882813 C 3.105469 -2.273438 3.117188 -1.917969 3.144531 -1.816406 C 3.167969 -1.714844 3.226563 -1.628906 3.320313 -1.566406 C 3.410156 -1.496094 3.523438 -1.464844 3.65625 -1.46875 C 3.835938 -1.464844 4.097656 -1.527344 4.449219 -1.660156 L 4.621094 -0.125 C 4.15625 0.0703125 3.636719 0.164063 3.058594 0.167969 C 2.699219 0.164063 2.375 0.105469 2.09375 -0.0117188 C 1.804688 -0.128906 1.597656 -0.28125 1.464844 -0.472656 C 1.332031 -0.660156 1.238281 -0.917969 1.1875 -1.246094 C 1.144531 -1.472656 1.125 -1.9375 1.125 -2.636719 L 1.125 -5.890625 L 0.21875 -5.890625 L 0.21875 -7.46875 L 1.125 -7.46875 L 1.125 -8.949219 L 3.109375 -10.105469 L 3.109375 -7.46875 Z M 4.457031 -7.46875 "/>
</symbol>
<symbol overflow="visible" id="glyph1-5">
<path style="stroke:none;" d="M 2.925781 0 L 0.949219 0 L 0.949219 -7.46875 L 2.785156 -7.46875 L 2.785156 -6.40625 C 3.09375 -6.902344 3.375 -7.234375 3.628906 -7.394531 C 3.878906 -7.554688 4.164063 -7.632813 4.484375 -7.636719 C 4.929688 -7.632813 5.363281 -7.507813 5.785156 -7.261719 L 5.175781 -5.539063 C 4.839844 -5.75 4.53125 -5.859375 4.246094 -5.863281 C 3.96875 -5.859375 3.734375 -5.78125 3.542969 -5.632813 C 3.347656 -5.476563 3.195313 -5.203125 3.089844 -4.808594 C 2.976563 -4.40625 2.921875 -3.570313 2.925781 -2.304688 Z M 2.925781 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-6">
<path style="stroke:none;" d="M 0.949219 0 L 0.949219 -10.308594 L 2.925781 -10.308594 L 2.925781 -6.59375 C 3.53125 -7.285156 4.253906 -7.632813 5.089844 -7.636719 C 5.996094 -7.632813 6.75 -7.304688 7.347656 -6.648438 C 7.941406 -5.988281 8.238281 -5.042969 8.242188 -3.8125 C 8.238281 -2.535156 7.933594 -1.550781 7.328125 -0.863281 C 6.71875 -0.175781 5.980469 0.164063 5.117188 0.167969 C 4.6875 0.164063 4.269531 0.0585938 3.855469 -0.152344 C 3.441406 -0.363281 3.082031 -0.675781 2.785156 -1.097656 L 2.785156 0 Z M 2.910156 -3.894531 C 2.90625 -3.117188 3.027344 -2.546875 3.277344 -2.179688 C 3.613281 -1.652344 4.070313 -1.386719 4.640625 -1.390625 C 5.074219 -1.386719 5.445313 -1.574219 5.753906 -1.949219 C 6.058594 -2.320313 6.210938 -2.90625 6.214844 -3.710938 C 6.210938 -4.5625 6.054688 -5.179688 5.75 -5.558594 C 5.4375 -5.933594 5.042969 -6.121094 4.5625 -6.125 C 4.085938 -6.121094 3.691406 -5.9375 3.378906 -5.570313 C 3.0625 -5.199219 2.90625 -4.640625 2.910156 -3.894531 Z M 2.910156 -3.894531 "/>
</symbol>
<symbol overflow="visible" id="glyph1-7">
<path style="stroke:none;" d="M 5.949219 0 L 5.949219 -1.117188 C 5.671875 -0.714844 5.316406 -0.402344 4.875 -0.175781 C 4.429688 0.0507813 3.960938 0.164063 3.472656 0.167969 C 2.96875 0.164063 2.519531 0.0585938 2.125 -0.160156 C 1.722656 -0.378906 1.433594 -0.691406 1.257813 -1.089844 C 1.078125 -1.488281 0.988281 -2.039063 0.992188 -2.742188 L 0.992188 -7.46875 L 2.96875 -7.46875 L 2.96875 -4.035156 C 2.964844 -2.984375 3 -2.339844 3.074219 -2.105469 C 3.144531 -1.863281 3.277344 -1.675781 3.472656 -1.542969 C 3.664063 -1.402344 3.90625 -1.335938 4.203125 -1.335938 C 4.539063 -1.335938 4.84375 -1.425781 5.109375 -1.613281 C 5.375 -1.792969 5.558594 -2.023438 5.660156 -2.300781 C 5.757813 -2.574219 5.804688 -3.246094 5.808594 -4.316406 L 5.808594 -7.46875 L 7.785156 -7.46875 L 7.785156 0 Z M 5.949219 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-8">
<path style="stroke:none;" d="M 0.578125 -3.839844 C 0.574219 -4.492188 0.734375 -5.128906 1.0625 -5.742188 C 1.382813 -6.355469 1.839844 -6.824219 2.433594 -7.148438 C 3.023438 -7.472656 3.6875 -7.632813 4.421875 -7.636719 C 5.550781 -7.632813 6.476563 -7.265625 7.199219 -6.535156 C 7.917969 -5.796875 8.277344 -4.871094 8.28125 -3.753906 C 8.277344 -2.621094 7.914063 -1.683594 7.1875 -0.945313 C 6.457031 -0.203125 5.539063 0.164063 4.4375 0.167969 C 3.75 0.164063 3.097656 0.0117188 2.476563 -0.292969 C 1.855469 -0.601563 1.382813 -1.054688 1.0625 -1.652344 C 0.734375 -2.25 0.574219 -2.976563 0.578125 -3.839844 Z M 2.601563 -3.734375 C 2.601563 -2.988281 2.777344 -2.421875 3.128906 -2.03125 C 3.480469 -1.636719 3.914063 -1.441406 4.429688 -1.441406 C 4.945313 -1.441406 5.375 -1.636719 5.726563 -2.03125 C 6.070313 -2.421875 6.246094 -2.992188 6.25 -3.746094 C 6.246094 -4.472656 6.070313 -5.035156 5.726563 -5.433594 C 5.375 -5.824219 4.945313 -6.023438 4.429688 -6.027344 C 3.914063 -6.023438 3.480469 -5.824219 3.128906 -5.433594 C 2.777344 -5.035156 2.601563 -4.46875 2.601563 -3.734375 Z M 2.601563 -3.734375 "/>
</symbol>
<symbol overflow="visible" id="glyph1-9">
<path style="stroke:none;" d="M 7.824219 0 L 5.851563 0 L 5.851563 -3.8125 C 5.847656 -4.613281 5.804688 -5.132813 5.722656 -5.375 C 5.636719 -5.609375 5.5 -5.792969 5.3125 -5.925781 C 5.121094 -6.054688 4.890625 -6.121094 4.625 -6.125 C 4.28125 -6.121094 3.976563 -6.027344 3.703125 -5.84375 C 3.429688 -5.652344 3.242188 -5.40625 3.144531 -5.097656 C 3.042969 -4.785156 2.992188 -4.210938 2.996094 -3.382813 L 2.996094 0 L 1.019531 0 L 1.019531 -7.46875 L 2.855469 -7.46875 L 2.855469 -6.371094 C 3.503906 -7.210938 4.324219 -7.632813 5.316406 -7.636719 C 5.746094 -7.632813 6.144531 -7.554688 6.507813 -7.398438 C 6.867188 -7.238281 7.140625 -7.039063 7.328125 -6.796875 C 7.511719 -6.554688 7.640625 -6.277344 7.714844 -5.96875 C 7.785156 -5.65625 7.820313 -5.214844 7.824219 -4.640625 Z M 7.824219 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-10">
<path style="stroke:none;" d=""/>
</symbol>
<symbol overflow="visible" id="glyph1-11">
<path style="stroke:none;" d="M 0.167969 -7.46875 L 1.265625 -7.46875 L 1.265625 -8.03125 C 1.265625 -8.65625 1.332031 -9.125 1.464844 -9.433594 C 1.597656 -9.742188 1.84375 -9.992188 2.203125 -10.191406 C 2.5625 -10.382813 3.015625 -10.480469 3.566406 -10.484375 C 4.125 -10.480469 4.675781 -10.398438 5.21875 -10.230469 L 4.949219 -8.851563 C 4.632813 -8.925781 4.332031 -8.964844 4.042969 -8.964844 C 3.753906 -8.964844 3.546875 -8.894531 3.425781 -8.761719 C 3.300781 -8.625 3.238281 -8.371094 3.242188 -7.996094 L 3.242188 -7.46875 L 4.71875 -7.46875 L 4.71875 -5.914063 L 3.242188 -5.914063 L 3.242188 0 L 1.265625 0 L 1.265625 -5.914063 L 0.167969 -5.914063 Z M 0.167969 -7.46875 "/>
</symbol>
<symbol overflow="visible" id="glyph1-12">
<path style="stroke:none;" d="M 3.367188 0 L 3.367188 -8.5625 L 0.308594 -8.5625 L 0.308594 -10.308594 L 8.5 -10.308594 L 8.5 -8.5625 L 5.449219 -8.5625 L 5.449219 0 Z M 3.367188 0 "/>
</symbol>
<symbol overflow="visible" id="glyph1-13">
<path style="stroke:none;" d="M 0.0976563 -7.46875 L 2.199219 -7.46875 L 3.988281 -2.164063 L 5.730469 -7.46875 L 7.777344 -7.46875 L 5.140625 -0.28125 L 4.667969 1.019531 C 4.492188 1.453125 4.328125 1.785156 4.171875 2.015625 C 4.015625 2.246094 3.832031 2.433594 3.628906 2.578125 C 3.421875 2.71875 3.171875 2.828125 2.878906 2.910156 C 2.578125 2.988281 2.242188 3.027344 1.871094 3.03125 C 1.488281 3.027344 1.117188 2.988281 0.753906 2.910156 L 0.578125 1.363281 C 0.882813 1.421875 1.160156 1.453125 1.414063 1.457031 C 1.867188 1.453125 2.207031 1.316406 2.429688 1.050781 C 2.648438 0.777344 2.816406 0.433594 2.9375 0.0195313 Z M 0.0976563 -7.46875 "/>
</symbol>
<symbol overflow="visible" id="glyph1-14">
<path style="stroke:none;" d="M 0.976563 -7.46875 L 2.820313 -7.46875 L 2.820313 -6.371094 C 3.054688 -6.742188 3.378906 -7.046875 3.789063 -7.285156 C 4.195313 -7.515625 4.648438 -7.632813 5.148438 -7.636719 C 6.011719 -7.632813 6.746094 -7.292969 7.355469 -6.617188 C 7.957031 -5.933594 8.261719 -4.988281 8.261719 -3.777344 C 8.261719 -2.527344 7.957031 -1.558594 7.347656 -0.867188 C 6.738281 -0.179688 6 0.164063 5.132813 0.167969 C 4.71875 0.164063 4.34375 0.0859375 4.011719 -0.078125 C 3.671875 -0.238281 3.320313 -0.519531 2.953125 -0.921875 L 2.953125 2.839844 L 0.976563 2.839844 Z M 2.933594 -3.859375 C 2.929688 -3.019531 3.09375 -2.398438 3.429688 -2 C 3.757813 -1.59375 4.164063 -1.394531 4.648438 -1.398438 C 5.101563 -1.394531 5.484375 -1.578125 5.792969 -1.949219 C 6.09375 -2.316406 6.246094 -2.921875 6.25 -3.761719 C 6.246094 -4.542969 6.089844 -5.121094 5.777344 -5.503906 C 5.464844 -5.878906 5.074219 -6.070313 4.613281 -6.074219 C 4.125 -6.070313 3.726563 -5.882813 3.410156 -5.515625 C 3.089844 -5.140625 2.929688 -4.589844 2.933594 -3.859375 Z M 2.933594 -3.859375 "/>
</symbol>
<symbol overflow="visible" id="glyph1-15">
<path style="stroke:none;" d="M 5.359375 -2.375 L 7.328125 -2.046875 C 7.070313 -1.320313 6.667969 -0.773438 6.125 -0.398438 C 5.578125 -0.0234375 4.898438 0.164063 4.078125 0.167969 C 2.777344 0.164063 1.816406 -0.257813 1.195313 -1.105469 C 0.703125 -1.78125 0.457031 -2.636719 0.457031 -3.675781 C 0.457031 -4.910156 0.777344 -5.882813 1.425781 -6.585938 C 2.070313 -7.285156 2.890625 -7.632813 3.882813 -7.636719 C 4.988281 -7.632813 5.863281 -7.265625 6.507813 -6.535156 C 7.148438 -5.796875 7.457031 -4.675781 7.433594 -3.164063 L 2.480469 -3.164063 C 2.492188 -2.578125 2.652344 -2.121094 2.960938 -1.796875 C 3.261719 -1.46875 3.640625 -1.304688 4.097656 -1.308594 C 4.402344 -1.304688 4.664063 -1.390625 4.878906 -1.558594 C 5.085938 -1.726563 5.246094 -1.996094 5.359375 -2.375 Z M 5.46875 -4.375 C 5.453125 -4.941406 5.308594 -5.375 5.027344 -5.675781 C 4.746094 -5.972656 4.402344 -6.121094 4 -6.125 C 3.566406 -6.121094 3.210938 -5.964844 2.933594 -5.652344 C 2.648438 -5.335938 2.507813 -4.910156 2.515625 -4.375 Z M 5.46875 -4.375 "/>
</symbol>
<symbol overflow="visible" id="glyph1-16">
<path style="stroke:none;" d="M 0.625 -5.089844 C 0.621094 -6.136719 0.777344 -7.019531 1.097656 -7.734375 C 1.328125 -8.257813 1.648438 -8.726563 2.054688 -9.148438 C 2.457031 -9.5625 2.902344 -9.871094 3.390625 -10.074219 C 4.027344 -10.34375 4.765625 -10.480469 5.609375 -10.484375 C 7.125 -10.480469 8.34375 -10.011719 9.257813 -9.070313 C 10.167969 -8.125 10.621094 -6.8125 10.625 -5.140625 C 10.621094 -3.472656 10.167969 -2.171875 9.265625 -1.234375 C 8.359375 -0.292969 7.152344 0.175781 5.640625 0.175781 C 4.105469 0.175781 2.886719 -0.289063 1.980469 -1.226563 C 1.074219 -2.15625 0.621094 -3.445313 0.625 -5.089844 Z M 2.769531 -5.160156 C 2.765625 -3.992188 3.035156 -3.105469 3.578125 -2.503906 C 4.113281 -1.898438 4.796875 -1.597656 5.632813 -1.601563 C 6.457031 -1.597656 7.136719 -1.898438 7.671875 -2.496094 C 8.203125 -3.09375 8.472656 -3.988281 8.472656 -5.1875 C 8.472656 -6.367188 8.210938 -7.25 7.695313 -7.832031 C 7.171875 -8.410156 6.484375 -8.699219 5.632813 -8.703125 C 4.769531 -8.699219 4.078125 -8.40625 3.554688 -7.820313 C 3.027344 -7.230469 2.765625 -6.34375 2.769531 -5.160156 Z M 2.769531 -5.160156 "/>
</symbol>
<symbol overflow="visible" id="glyph1-17">
<path style="stroke:none;" d="M 2.511719 -5.1875 L 0.71875 -5.511719 C 0.917969 -6.230469 1.265625 -6.765625 1.757813 -7.113281 C 2.25 -7.460938 2.980469 -7.632813 3.953125 -7.636719 C 4.832031 -7.632813 5.488281 -7.53125 5.917969 -7.324219 C 6.347656 -7.113281 6.648438 -6.847656 6.828125 -6.527344 C 7 -6.207031 7.089844 -5.617188 7.09375 -4.761719 L 7.074219 -2.453125 C 7.070313 -1.792969 7.101563 -1.308594 7.167969 -1 C 7.226563 -0.6875 7.347656 -0.355469 7.523438 0 L 5.570313 0 C 5.515625 -0.128906 5.453125 -0.320313 5.378906 -0.582031 C 5.34375 -0.695313 5.320313 -0.773438 5.308594 -0.816406 C 4.96875 -0.484375 4.605469 -0.238281 4.222656 -0.078125 C 3.835938 0.0859375 3.425781 0.164063 2.996094 0.167969 C 2.222656 0.164063 1.617188 -0.0429688 1.175781 -0.457031 C 0.730469 -0.871094 0.507813 -1.398438 0.511719 -2.039063 C 0.507813 -2.460938 0.609375 -2.835938 0.8125 -3.167969 C 1.011719 -3.496094 1.292969 -3.75 1.660156 -3.925781 C 2.019531 -4.101563 2.546875 -4.253906 3.234375 -4.386719 C 4.15625 -4.558594 4.792969 -4.71875 5.152344 -4.871094 L 5.152344 -5.070313 C 5.148438 -5.445313 5.054688 -5.71875 4.871094 -5.882813 C 4.679688 -6.042969 4.328125 -6.121094 3.8125 -6.125 C 3.457031 -6.121094 3.183594 -6.054688 2.988281 -5.917969 C 2.789063 -5.777344 2.628906 -5.53125 2.511719 -5.1875 Z M 5.152344 -3.585938 C 4.894531 -3.5 4.496094 -3.398438 3.949219 -3.285156 C 3.402344 -3.164063 3.042969 -3.046875 2.875 -2.9375 C 2.613281 -2.75 2.484375 -2.519531 2.488281 -2.242188 C 2.484375 -1.964844 2.585938 -1.726563 2.796875 -1.523438 C 3 -1.320313 3.265625 -1.21875 3.585938 -1.222656 C 3.941406 -1.21875 4.28125 -1.335938 4.605469 -1.574219 C 4.84375 -1.75 5 -1.96875 5.078125 -2.230469 C 5.125 -2.394531 5.148438 -2.714844 5.152344 -3.191406 Z M 5.152344 -3.585938 "/>
</symbol>
<symbol overflow="visible" id="glyph2-0">
<path style="stroke:none;" d="M 1.199219 0 L 1.199219 -6 L 6 -6 L 6 0 Z M 1.351563 -0.148438 L 5.851563 -0.148438 L 5.851563 -5.851563 L 1.351563 -5.851563 Z M 1.351563 -0.148438 "/>
</symbol>
<symbol overflow="visible" id="glyph2-1">
<path style="stroke:none;" d="M 5.644531 -2.410156 L 6.554688 -2.179688 C 6.359375 -1.429688 6.015625 -0.859375 5.523438 -0.46875 C 5.027344 -0.078125 4.421875 0.117188 3.707031 0.117188 C 2.964844 0.117188 2.363281 -0.03125 1.898438 -0.335938 C 1.433594 -0.632813 1.078125 -1.070313 0.839844 -1.644531 C 0.59375 -2.214844 0.472656 -2.828125 0.476563 -3.488281 C 0.472656 -4.199219 0.609375 -4.824219 0.886719 -5.359375 C 1.15625 -5.890625 1.546875 -6.296875 2.054688 -6.574219 C 2.558594 -6.847656 3.113281 -6.984375 3.722656 -6.988281 C 4.40625 -6.984375 4.984375 -6.808594 5.457031 -6.460938 C 5.921875 -6.109375 6.25 -5.617188 6.4375 -4.988281 L 5.539063 -4.777344 C 5.375 -5.273438 5.144531 -5.636719 4.84375 -5.867188 C 4.539063 -6.09375 4.160156 -6.210938 3.703125 -6.210938 C 3.171875 -6.210938 2.730469 -6.082031 2.378906 -5.832031 C 2.023438 -5.574219 1.773438 -5.234375 1.628906 -4.8125 C 1.484375 -4.382813 1.410156 -3.945313 1.414063 -3.492188 C 1.410156 -2.90625 1.496094 -2.394531 1.667969 -1.960938 C 1.835938 -1.523438 2.101563 -1.199219 2.464844 -0.984375 C 2.820313 -0.765625 3.210938 -0.65625 3.632813 -0.660156 C 4.140625 -0.65625 4.570313 -0.804688 4.925781 -1.101563 C 5.277344 -1.394531 5.515625 -1.828125 5.644531 -2.410156 Z M 5.644531 -2.410156 "/>
</symbol>
<symbol overflow="visible" id="glyph2-2">
<path style="stroke:none;" d="M 2.488281 0 L 2.488281 -6.0625 L 0.226563 -6.0625 L 0.226563 -6.871094 L 5.671875 -6.871094 L 5.671875 -6.0625 L 3.398438 -6.0625 L 3.398438 0 Z M 2.488281 0 "/>
</symbol>
<symbol overflow="visible" id="glyph2-3">
<path style="stroke:none;" d="M 0.753906 0 L 0.753906 -6.871094 L 3.800781 -6.871094 C 4.410156 -6.867188 4.875 -6.804688 5.195313 -6.683594 C 5.511719 -6.558594 5.765625 -6.339844 5.960938 -6.03125 C 6.148438 -5.714844 6.246094 -5.371094 6.25 -4.996094 C 6.246094 -4.507813 6.085938 -4.097656 5.773438 -3.761719 C 5.453125 -3.425781 4.96875 -3.210938 4.3125 -3.125 C 4.550781 -3.007813 4.730469 -2.894531 4.859375 -2.785156 C 5.121094 -2.535156 5.375 -2.230469 5.617188 -1.871094 L 6.8125 0 L 5.667969 0 L 4.757813 -1.429688 C 4.492188 -1.839844 4.273438 -2.152344 4.101563 -2.375 C 3.929688 -2.589844 3.773438 -2.746094 3.640625 -2.835938 C 3.5 -2.921875 3.363281 -2.980469 3.226563 -3.019531 C 3.121094 -3.035156 2.953125 -3.046875 2.71875 -3.050781 L 1.664063 -3.050781 L 1.664063 0 Z M 1.664063 -3.839844 L 3.617188 -3.839844 C 4.03125 -3.835938 4.359375 -3.878906 4.59375 -3.96875 C 4.828125 -4.050781 5.003906 -4.1875 5.128906 -4.378906 C 5.246094 -4.566406 5.308594 -4.773438 5.3125 -4.996094 C 5.308594 -5.320313 5.191406 -5.585938 4.957031 -5.796875 C 4.71875 -6.003906 4.34375 -6.109375 3.839844 -6.113281 L 1.664063 -6.113281 Z M 1.664063 -3.839844 "/>
</symbol>
<symbol overflow="visible" id="glyph2-4">
<path style="stroke:none;" d="M 0.703125 0 L 0.703125 -6.871094 L 1.613281 -6.871094 L 1.613281 -0.8125 L 4.996094 -0.8125 L 4.996094 0 Z M 0.703125 0 "/>
</symbol>
<symbol overflow="visible" id="glyph2-5">
<path style="stroke:none;" d="M 0.851563 -4.015625 L 0.851563 -4.976563 L 1.8125 -4.976563 L 1.8125 -4.015625 Z M 0.851563 0 L 0.851563 -0.960938 L 1.8125 -0.960938 L 1.8125 0 C 1.808594 0.351563 1.746094 0.636719 1.625 0.855469 C 1.496094 1.070313 1.300781 1.238281 1.03125 1.359375 L 0.796875 1 C 0.972656 0.917969 1.101563 0.800781 1.1875 0.652344 C 1.269531 0.496094 1.316406 0.28125 1.332031 0 Z M 0.851563 0 "/>
</symbol>
<symbol overflow="visible" id="glyph2-6">
<path style="stroke:none;" d="M 0.757813 0 L 0.757813 -6.871094 L 5.726563 -6.871094 L 5.726563 -6.0625 L 1.667969 -6.0625 L 1.667969 -3.957031 L 5.46875 -3.957031 L 5.46875 -3.148438 L 1.667969 -3.148438 L 1.667969 -0.8125 L 5.886719 -0.8125 L 5.886719 0 Z M 0.757813 0 "/>
</symbol>
<symbol overflow="visible" id="glyph2-7">
<path style="stroke:none;" d="M 0.0429688 0 L 2.699219 -3.582031 L 0.355469 -6.871094 L 1.4375 -6.871094 L 2.6875 -5.109375 C 2.941406 -4.742188 3.125 -4.460938 3.238281 -4.265625 C 3.390625 -4.515625 3.570313 -4.773438 3.78125 -5.046875 L 5.164063 -6.871094 L 6.15625 -6.871094 L 3.742188 -3.632813 L 6.34375 0 L 5.21875 0 L 3.488281 -2.453125 C 3.386719 -2.589844 3.289063 -2.742188 3.1875 -2.910156 C 3.03125 -2.65625 2.921875 -2.484375 2.859375 -2.394531 L 1.132813 0 Z M 0.0429688 0 "/>
</symbol>
<symbol overflow="visible" id="glyph2-8">
<path style="stroke:none;" d="M 0.742188 0 L 0.742188 -6.871094 L 3.109375 -6.871094 C 3.640625 -6.867188 4.046875 -6.835938 4.332031 -6.773438 C 4.722656 -6.679688 5.058594 -6.515625 5.339844 -6.28125 C 5.699219 -5.972656 5.972656 -5.578125 6.152344 -5.105469 C 6.332031 -4.625 6.421875 -4.082031 6.421875 -3.472656 C 6.421875 -2.949219 6.359375 -2.488281 6.238281 -2.085938 C 6.113281 -1.679688 5.957031 -1.34375 5.769531 -1.082031 C 5.578125 -0.816406 5.371094 -0.609375 5.144531 -0.460938 C 4.917969 -0.308594 4.644531 -0.195313 4.324219 -0.117188 C 4.003906 -0.0390625 3.632813 0 3.21875 0 Z M 1.648438 -0.8125 L 3.117188 -0.8125 C 3.570313 -0.808594 3.925781 -0.851563 4.183594 -0.9375 C 4.441406 -1.019531 4.644531 -1.136719 4.800781 -1.292969 C 5.011719 -1.507813 5.179688 -1.796875 5.304688 -2.164063 C 5.421875 -2.523438 5.484375 -2.964844 5.484375 -3.488281 C 5.484375 -4.203125 5.363281 -4.757813 5.128906 -5.144531 C 4.890625 -5.527344 4.605469 -5.785156 4.269531 -5.921875 C 4.023438 -6.011719 3.632813 -6.058594 3.09375 -6.0625 L 1.648438 -6.0625 Z M 1.648438 -0.8125 "/>
</symbol>
<symbol overflow="visible" id="glyph2-9">
<path style="stroke:none;" d="M 0.710938 0 L 0.710938 -6.871094 L 2.082031 -6.871094 L 3.707031 -2.007813 C 3.855469 -1.550781 3.964844 -1.210938 4.035156 -0.988281 C 4.109375 -1.234375 4.230469 -1.601563 4.402344 -2.089844 L 6.046875 -6.871094 L 7.269531 -6.871094 L 7.269531 0 L 6.394531 0 L 6.394531 -5.75 L 4.398438 0 L 3.578125 0 L 1.589844 -5.851563 L 1.589844 0 Z M 0.710938 0 "/>
</symbol>
<symbol overflow="visible" id="glyph2-10">
<path style="stroke:none;" d="M 0.894531 0 L 0.894531 -6.871094 L 1.804688 -6.871094 L 1.804688 0 Z M 0.894531 0 "/>
</symbol>
<symbol overflow="visible" id="glyph2-11">
<path style="stroke:none;" d="M 0.730469 0 L 0.730469 -6.871094 L 1.664063 -6.871094 L 5.273438 -1.476563 L 5.273438 -6.871094 L 6.144531 -6.871094 L 6.144531 0 L 5.210938 0 L 1.601563 -5.398438 L 1.601563 0 Z M 0.730469 0 "/>
</symbol>
</g>
<clipPath id="clip1">
  <path d="M 207 59.039063 L 330 59.039063 L 330 106 L 207 106 Z M 207 59.039063 "/>
</clipPath>
<clipPath id="clip2">
  <path d="M 207 59.039063 L 330.757813 59.039063 L 330.757813 106 L 207 106 Z M 207 59.039063 "/>
</clipPath>
</defs>
<g id="surface28">
<rect x="0" y="0" width="360" height="360" style="fill:rgb(100%,100%,100%);fill-opacity:1;stroke:none;"/>
<path style="fill-rule:nonzero;fill:rgb(20%,13.333333%,53.333333%);fill-opacity:1;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 278.667969 172.800781 L 278.625 170.097656 L 278.492188 167.402344 L 278.277344 164.707031 L 277.976563 162.023438 L 277.585938 159.351563 L 277.113281 156.691406 L 276.554688 154.050781 L 275.910156 151.425781 L 275.183594 148.824219 L 274.375 146.246094 L 273.480469 143.695313 L 272.507813 141.175781 L 271.453125 138.691406 L 270.320313 136.238281 L 269.109375 133.824219 L 267.824219 131.449219 L 266.460938 129.117188 L 265.023438 126.828125 L 263.511719 124.589844 L 261.933594 122.398438 L 260.28125 120.261719 L 258.566406 118.175781 L 256.78125 116.148438 L 254.933594 114.175781 L 253.023438 112.265625 L 251.050781 110.417969 L 249.023438 108.636719 L 246.9375 106.917969 L 244.800781 105.265625 L 242.609375 103.6875 L 240.371094 102.175781 L 238.082031 100.738281 L 235.75 99.375 L 233.375 98.089844 L 230.960938 96.878906 L 228.507813 95.746094 L 226.023438 94.691406 L 223.503906 93.71875 L 220.953125 92.828125 L 218.375 92.015625 L 215.773438 91.289063 L 213.152344 90.644531 L 210.507813 90.085938 L 207.847656 89.613281 L 205.175781 89.226563 L 202.492188 88.921875 L 199.800781 88.707031 L 197.101563 88.578125 L 194.398438 88.535156 L 194.398438 172.800781 Z M 278.667969 172.800781 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 253.984375 113.214844 L 256.964844 110.234375 "/>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph0-1" x="259.945313" y="111.464844"/>
  <use xlink:href="#glyph0-2" x="266.619141" y="111.464844"/>
  <use xlink:href="#glyph0-3" x="273.292969" y="111.464844"/>
</g>
<path style="fill-rule:nonzero;fill:rgb(53.333333%,80%,93.333333%);fill-opacity:1;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 194.398438 88.535156 L 191.699219 88.578125 L 189 88.707031 L 186.308594 88.921875 L 183.625 89.226563 L 180.949219 89.613281 L 178.292969 90.085938 L 175.648438 90.644531 L 173.023438 91.289063 L 170.421875 92.015625 L 167.847656 92.828125 L 165.296875 93.71875 L 162.777344 94.691406 L 160.289063 95.746094 L 157.839844 96.878906 L 155.421875 98.089844 L 153.050781 99.375 L 150.714844 100.738281 L 148.429688 102.175781 L 146.191406 103.6875 L 144 105.265625 L 141.859375 106.917969 L 139.777344 108.636719 L 137.746094 110.417969 L 135.777344 112.265625 L 133.867188 114.175781 L 132.019531 116.148438 L 130.234375 118.175781 L 128.519531 120.261719 L 126.867188 122.398438 L 125.285156 124.589844 L 123.777344 126.828125 L 122.339844 129.117188 L 120.976563 131.449219 L 119.6875 133.824219 L 118.476563 136.238281 L 117.34375 138.691406 L 116.292969 141.175781 L 115.320313 143.695313 L 114.425781 146.246094 L 113.617188 148.824219 L 112.890625 151.425781 L 112.246094 154.050781 L 111.6875 156.691406 L 111.214844 159.351563 L 110.824219 162.023438 L 110.523438 164.707031 L 110.304688 167.402344 L 110.175781 170.097656 L 110.132813 172.800781 L 194.398438 172.800781 Z M 194.398438 88.535156 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 134.816406 113.214844 L 131.835938 110.234375 "/>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph0-1" x="104.839844" y="111.464844"/>
  <use xlink:href="#glyph0-2" x="111.513672" y="111.464844"/>
  <use xlink:href="#glyph0-3" x="118.1875" y="111.464844"/>
</g>
<path style="fill-rule:nonzero;fill:rgb(26.666667%,66.666667%,60%);fill-opacity:1;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 110.132813 172.800781 L 110.175781 175.472656 L 110.304688 178.144531 L 110.515625 180.808594 L 110.8125 183.46875 L 111.191406 186.113281 L 111.65625 188.746094 L 112.203125 191.363281 L 112.835938 193.964844 L 113.546875 196.539063 L 114.339844 199.09375 L 115.214844 201.621094 L 116.167969 204.117188 L 117.203125 206.585938 L 118.3125 209.015625 L 119.5 211.414063 L 120.761719 213.769531 L 122.101563 216.085938 L 123.511719 218.359375 L 124.992188 220.585938 L 126.542969 222.761719 L 128.160156 224.890625 L 129.847656 226.964844 L 131.597656 228.988281 L 133.414063 230.949219 L 135.289063 232.855469 L 137.222656 234.703125 L 139.21875 236.484375 L 141.265625 238.203125 L 143.367188 239.855469 L 145.519531 241.441406 L 147.722656 242.957031 L 149.972656 244.402344 L 152.265625 245.777344 L 154.601563 247.078125 L 156.980469 248.300781 L 159.394531 249.453125 L 161.84375 250.523438 L 164.328125 251.515625 L 166.839844 252.433594 L 169.378906 253.265625 L 171.945313 254.019531 L 174.535156 254.691406 L 177.140625 255.28125 L 179.765625 255.785156 L 182.40625 256.207031 L 185.058594 256.546875 L 187.722656 256.800781 L 190.390625 256.972656 L 193.0625 257.054688 L 195.738281 257.054688 L 198.410156 256.972656 L 201.078125 256.800781 L 203.738281 256.546875 L 206.390625 256.207031 L 209.03125 255.785156 L 211.660156 255.28125 L 214.265625 254.691406 L 216.855469 254.019531 L 219.421875 253.265625 L 221.960938 252.433594 L 224.472656 251.515625 L 226.957031 250.523438 L 229.40625 249.453125 L 231.820313 248.300781 L 234.195313 247.078125 L 236.535156 245.777344 L 238.828125 244.402344 L 241.078125 242.957031 L 243.28125 241.441406 L 245.433594 239.855469 L 247.535156 238.203125 L 249.582031 236.484375 L 251.574219 234.703125 L 253.511719 232.855469 L 255.386719 230.949219 L 257.199219 228.988281 L 258.953125 226.964844 L 260.636719 224.890625 L 262.257813 222.761719 L 263.808594 220.585938 L 265.289063 218.359375 L 266.699219 216.085938 L 268.035156 213.769531 L 269.300781 211.414063 L 270.488281 209.015625 L 271.597656 206.585938 L 272.628906 204.117188 L 273.585938 201.621094 L 274.460938 199.09375 L 275.253906 196.539063 L 275.964844 193.964844 L 276.597656 191.363281 L 277.144531 188.746094 L 277.609375 186.113281 L 277.988281 183.46875 L 278.285156 180.808594 L 278.496094 178.144531 L 278.625 175.472656 L 278.667969 172.800781 Z M 110.132813 172.800781 "/>
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 194.398438 257.066406 L 194.398438 261.28125 "/>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph0-2" x="170.382813" y="269.703125"/>
  <use xlink:href="#glyph0-4" x="177.056641" y="269.703125"/>
  <use xlink:href="#glyph0-3" x="183.730469" y="269.703125"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph1-1" x="73.59375" y="34.675781"/>
  <use xlink:href="#glyph1-2" x="83.992969" y="34.675781"/>
  <use xlink:href="#glyph1-3" x="87.99375" y="34.675781"/>
  <use xlink:href="#glyph1-4" x="96.002344" y="34.675781"/>
  <use xlink:href="#glyph1-5" x="100.797656" y="34.675781"/>
  <use xlink:href="#glyph1-2" x="106.401563" y="34.675781"/>
  <use xlink:href="#glyph1-6" x="110.402344" y="34.675781"/>
  <use xlink:href="#glyph1-7" x="119.198438" y="34.675781"/>
  <use xlink:href="#glyph1-4" x="127.994531" y="34.675781"/>
  <use xlink:href="#glyph1-2" x="132.789844" y="34.675781"/>
  <use xlink:href="#glyph1-8" x="136.790625" y="34.675781"/>
  <use xlink:href="#glyph1-9" x="145.586719" y="34.675781"/>
  <use xlink:href="#glyph1-10" x="154.382813" y="34.675781"/>
  <use xlink:href="#glyph1-8" x="158.383594" y="34.675781"/>
  <use xlink:href="#glyph1-11" x="167.179688" y="34.675781"/>
  <use xlink:href="#glyph1-10" x="171.975" y="34.675781"/>
  <use xlink:href="#glyph1-12" x="175.975781" y="34.675781"/>
  <use xlink:href="#glyph1-13" x="184.771875" y="34.675781"/>
  <use xlink:href="#glyph1-14" x="192.780469" y="34.675781"/>
  <use xlink:href="#glyph1-15" x="201.576562" y="34.675781"/>
  <use xlink:href="#glyph1-3" x="209.585156" y="34.675781"/>
  <use xlink:href="#glyph1-10" x="217.59375" y="34.675781"/>
  <use xlink:href="#glyph1-8" x="221.594531" y="34.675781"/>
  <use xlink:href="#glyph1-11" x="230.390625" y="34.675781"/>
  <use xlink:href="#glyph1-10" x="235.185937" y="34.675781"/>
  <use xlink:href="#glyph1-16" x="239.186719" y="34.675781"/>
  <use xlink:href="#glyph1-14" x="250.3875" y="34.675781"/>
  <use xlink:href="#glyph1-15" x="259.183594" y="34.675781"/>
  <use xlink:href="#glyph1-5" x="267.192187" y="34.675781"/>
  <use xlink:href="#glyph1-17" x="272.796094" y="34.675781"/>
  <use xlink:href="#glyph1-4" x="280.804687" y="34.675781"/>
  <use xlink:href="#glyph1-2" x="285.6" y="34.675781"/>
  <use xlink:href="#glyph1-8" x="289.600781" y="34.675781"/>
  <use xlink:href="#glyph1-9" x="298.396875" y="34.675781"/>
  <use xlink:href="#glyph1-3" x="307.192969" y="34.675781"/>
</g>
<g clip-path="url(#clip1)" clip-rule="nonzero">
<path style=" stroke:none;fill-rule:nonzero;fill:rgb(100%,100%,100%);fill-opacity:1;" d="M 207.894531 59.039063 L 329.757813 59.039063 L 329.757813 105.117188 L 207.894531 105.117188 Z M 207.894531 59.039063 "/>
</g>
<g clip-path="url(#clip2)" clip-rule="nonzero">
<path style="fill:none;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 207.894531 59.039063 L 329.757813 59.039063 L 329.757813 105.117188 L 207.894531 105.117188 Z M 207.894531 59.039063 "/>
</g>
<path style="fill-rule:nonzero;fill:rgb(20%,13.333333%,53.333333%);fill-opacity:1;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 216.535156 67.679688 L 223.445313 67.679688 L 223.445313 73.441406 L 216.535156 73.441406 Z M 216.535156 67.679688 "/>
<path style="fill-rule:nonzero;fill:rgb(53.333333%,80%,93.333333%);fill-opacity:1;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 216.535156 79.199219 L 223.445313 79.199219 L 223.445313 84.960938 L 216.535156 84.960938 Z M 216.535156 79.199219 "/>
<path style="fill-rule:nonzero;fill:rgb(26.666667%,66.666667%,60%);fill-opacity:1;stroke-width:0.75;stroke-linecap:round;stroke-linejoin:round;stroke:rgb(0%,0%,0%);stroke-opacity:1;stroke-miterlimit:10;" d="M 216.535156 90.71875 L 223.445313 90.71875 L 223.445313 96.480469 L 216.535156 96.480469 Z M 216.535156 90.71875 "/>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-1" x="232.089844" y="73.996094"/>
  <use xlink:href="#glyph2-2" x="239.022656" y="73.996094"/>
  <use xlink:href="#glyph2-3" x="244.886719" y="73.996094"/>
  <use xlink:href="#glyph2-4" x="251.819531" y="73.996094"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-1" x="232.089844" y="85.515625"/>
  <use xlink:href="#glyph2-2" x="239.022656" y="85.515625"/>
  <use xlink:href="#glyph2-3" x="244.886719" y="85.515625"/>
  <use xlink:href="#glyph2-4" x="251.819531" y="85.515625"/>
  <use xlink:href="#glyph2-5" x="257.158594" y="85.515625"/>
  <use xlink:href="#glyph2-6" x="259.825781" y="85.515625"/>
  <use xlink:href="#glyph2-7" x="266.228906" y="85.515625"/>
  <use xlink:href="#glyph2-2" x="272.632031" y="85.515625"/>
  <use xlink:href="#glyph2-1" x="278.496094" y="85.515625"/>
  <use xlink:href="#glyph2-4" x="285.428906" y="85.515625"/>
  <use xlink:href="#glyph2-4" x="290.767969" y="85.515625"/>
  <use xlink:href="#glyph2-5" x="296.107031" y="85.515625"/>
  <use xlink:href="#glyph2-8" x="298.774219" y="85.515625"/>
  <use xlink:href="#glyph2-9" x="305.707031" y="85.515625"/>
  <use xlink:href="#glyph2-5" x="313.703906" y="85.515625"/>
  <use xlink:href="#glyph2-6" x="316.371094" y="85.515625"/>
  <use xlink:href="#glyph2-10" x="322.774219" y="85.515625"/>
</g>
<g style="fill:rgb(0%,0%,0%);fill-opacity:1;">
  <use xlink:href="#glyph2-1" x="232.089844" y="97.035156"/>
  <use xlink:href="#glyph2-2" x="239.022656" y="97.035156"/>
  <use xlink:href="#glyph2-3" x="244.886719" y="97.035156"/>
  <use xlink:href="#glyph2-4" x="251.819531" y="97.035156"/>
  <use xlink:href="#glyph2-5" x="257.158594" y="97.035156"/>
  <use xlink:href="#glyph2-6" x="259.825781" y="97.035156"/>
  <use xlink:href="#glyph2-7" x="266.228906" y="97.035156"/>
  <use xlink:href="#glyph2-2" x="272.632031" y="97.035156"/>
  <use xlink:href="#glyph2-1" x="278.496094" y="97.035156"/>
  <use xlink:href="#glyph2-4" x="285.428906" y="97.035156"/>
  <use xlink:href="#glyph2-4" x="290.767969" y="97.035156"/>
  <use xlink:href="#glyph2-5" x="296.107031" y="97.035156"/>
  <use xlink:href="#glyph2-10" x="298.774219" y="97.035156"/>
  <use xlink:href="#glyph2-11" x="301.441406" y="97.035156"/>
  <use xlink:href="#glyph2-2" x="308.374219" y="97.035156"/>
</g>
</g>
</svg>
